module alu (
  input  wire [31:0] a,
  input  wire [31:0] b,
  input  wire [3:0]  alu_ctrl,
  output reg  [31:0] result,
  output wire zero
);

assign zero = (result == 32'd0);

always @(*) begin
  result = 32'd0;
  case (alu_ctrl)
    4'b0000: result = a + b;               // ADD
    4'b0001: result = a - b;               // SUB
    4'b0010: result = a & b;               // AND
    4'b0011: result = a | b;               // OR
    4'b0100: result = (a < b) ? 32'd1 : 0; // SLT
    default: result = 32'd0;
  endcase
end

endmodule
