* NGSPICE file created from cpu_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

.subckt cpu_top VGND VPWR clk dbg_alu[0] dbg_alu[10] dbg_alu[11] dbg_alu[12] dbg_alu[13]
+ dbg_alu[14] dbg_alu[15] dbg_alu[16] dbg_alu[17] dbg_alu[18] dbg_alu[19] dbg_alu[1]
+ dbg_alu[20] dbg_alu[21] dbg_alu[22] dbg_alu[23] dbg_alu[24] dbg_alu[25] dbg_alu[26]
+ dbg_alu[27] dbg_alu[28] dbg_alu[29] dbg_alu[2] dbg_alu[30] dbg_alu[31] dbg_alu[3]
+ dbg_alu[4] dbg_alu[5] dbg_alu[6] dbg_alu[7] dbg_alu[8] dbg_alu[9] dbg_instr[0] dbg_instr[12]
+ dbg_instr[13] dbg_instr[14] dbg_instr[15] dbg_instr[16] dbg_instr[17] dbg_instr[18]
+ dbg_instr[19] dbg_instr[1] dbg_instr[20] dbg_instr[21] dbg_instr[22] dbg_instr[23]
+ dbg_instr[24] dbg_instr[25] dbg_instr[26] dbg_instr[27] dbg_instr[28] dbg_instr[2]
+ dbg_instr[30] dbg_instr[31] dbg_instr[3] dbg_instr[4] dbg_instr[5] dbg_mem_addr[0]
+ dbg_mem_addr[10] dbg_mem_addr[11] dbg_mem_addr[12] dbg_mem_addr[13] dbg_mem_addr[14]
+ dbg_mem_addr[15] dbg_mem_addr[16] dbg_mem_addr[17] dbg_mem_addr[18] dbg_mem_addr[19]
+ dbg_mem_addr[1] dbg_mem_addr[20] dbg_mem_addr[21] dbg_mem_addr[22] dbg_mem_addr[23]
+ dbg_mem_addr[24] dbg_mem_addr[25] dbg_mem_addr[26] dbg_mem_addr[27] dbg_mem_addr[28]
+ dbg_mem_addr[29] dbg_mem_addr[2] dbg_mem_addr[30] dbg_mem_addr[31] dbg_mem_addr[3]
+ dbg_mem_addr[4] dbg_mem_addr[5] dbg_mem_addr[6] dbg_mem_addr[7] dbg_mem_addr[8]
+ dbg_mem_addr[9] dbg_memread dbg_memwrite dbg_pc[10] dbg_pc[11] dbg_pc[12] dbg_pc[13]
+ dbg_pc[14] dbg_pc[15] dbg_pc[16] dbg_pc[17] dbg_pc[18] dbg_pc[19] dbg_pc[20] dbg_pc[21]
+ dbg_pc[22] dbg_pc[23] dbg_pc[24] dbg_pc[25] dbg_pc[26] dbg_pc[27] dbg_pc[28] dbg_pc[29]
+ dbg_pc[2] dbg_pc[30] dbg_pc[31] dbg_pc[3] dbg_pc[4] dbg_pc[5] dbg_pc[6] dbg_pc[7]
+ dbg_pc[8] dbg_pc[9] dbg_wb[0] dbg_wb[10] dbg_wb[11] dbg_wb[12] dbg_wb[13] dbg_wb[14]
+ dbg_wb[15] dbg_wb[16] dbg_wb[17] dbg_wb[18] dbg_wb[19] dbg_wb[1] dbg_wb[20] dbg_wb[21]
+ dbg_wb[22] dbg_wb[23] dbg_wb[24] dbg_wb[25] dbg_wb[26] dbg_wb[27] dbg_wb[28] dbg_wb[29]
+ dbg_wb[2] dbg_wb[30] dbg_wb[31] dbg_wb[3] dbg_wb[4] dbg_wb[5] dbg_wb[6] dbg_wb[7]
+ dbg_wb[8] dbg_wb[9] dbg_wb_rd[0] dbg_wb_rd[1] dbg_wb_rd[2] dbg_wb_rd[3] dbg_wb_we
+ rst dbg_instr[7] dbg_instr[6] dbg_pc[0] dbg_instr[29] dbg_instr[11] dbg_instr[10]
+ dbg_wb_rd[4] dbg_instr[9] dbg_instr[8] dbg_pc[1]
XFILLER_0_281_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2106_ _0766_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2037_ _0759_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__inv_2
XFILLER_0_210_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1064 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer7 _1003_ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__buf_2
XFILLER_0_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1270_ net80 net79 net78 _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__and4_2
XFILLER_0_78_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_283_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1606_ _0434_ _0435_ _0430_ _0431_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2586_ net31 VGND VGND VPWR VPWR _2586_/X sky130_fd_sc_hd__buf_2
XFILLER_0_125_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1537_ ID_EX.ex_rt_data\[10\] net197 VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1468_ _0954_ _1061_ _1062_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_199_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1399_ _0995_ _0997_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__xor2_2
XFILLER_0_241_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold170 net66 VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold181 RF.regs\[1\]\[26\] VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_258_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold192 net44 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2371_ clknet_leaf_25_clk net58 _0169_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1322_ _0935_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1253_ net269 _0897_ _0884_ _0898_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1184_ net288 _0865_ _0871_ _0868_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__a22o_1
XFILLER_0_194_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2569_ net118 VGND VGND VPWR VPWR _2569_/X sky130_fd_sc_hd__buf_2
XFILLER_0_273_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_242_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_528 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_9234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_9256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_267_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1940_ _0750_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1871_ _0315_ _0687_ _0634_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_910 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2354_ clknet_leaf_12_clk net213 _0152_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1305_ _0905_ _0924_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__and2b_1
XFILLER_0_276_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2285_ clknet_leaf_6_clk net300 _0083_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_263_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1236_ net233 _0895_ _0866_ _0894_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__a22o_1
XFILLER_0_237_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1167_ net239 _0853_ _0861_ _0855_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1098_ _0810_ MEM_WB.wb_alu_result\[19\] VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1036 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_259_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_284_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_266_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2070_ _0762_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1923_ _0704_ _0720_ _0736_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__and3_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1854_ _0573_ _0666_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_280_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_245_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1785_ net119 ID_EX.ex_rs_data\[23\] _0591_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2406_ clknet_leaf_0_clk _0303_ VGND VGND VPWR VPWR RF.regs\[1\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2337_ clknet_leaf_9_clk net25 _0135_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_224_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2268_ clknet_leaf_7_clk _0241_ _0066_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_240_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1219_ RF.regs\[1\]\[2\] _0849_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__and2_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2199_ _0748_ net125 _0773_ _0805_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__a31o_1
XFILLER_0_211_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold30 EX_MEM.mem_rd\[1\] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_264_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold41 ID_EX.ex_rt_data\[23\] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold52 _0234_ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold63 ID_EX.ex_rt_data\[16\] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold74 _0262_ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_242_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold85 ID_EX.ex_rt_data\[18\] VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_243_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold96 _0221_ VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_5 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_223_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1570_ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__buf_8
XFILLER_0_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2122_ _0767_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer17 _0321_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2053_ _0761_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__inv_2
Xrebuffer28 _1009_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1906_ _0704_ _0720_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1837_ _0383_ net59 _0573_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1768_ _0381_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__buf_4
XFILLER_0_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1699_ _0520_ _0521_ _0524_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__or3b_1
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_259_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput7 net7 VGND VGND VPWR VPWR dbg_alu[14] sky130_fd_sc_hd__clkbuf_4
Xoutput20 net20 VGND VGND VPWR VPWR dbg_alu[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput31 net31 VGND VGND VPWR VPWR dbg_alu[7] sky130_fd_sc_hd__buf_2
XFILLER_0_275_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput42 net42 VGND VGND VPWR VPWR dbg_mem_addr[10] sky130_fd_sc_hd__clkbuf_4
XTAP_6010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput53 net53 VGND VGND VPWR VPWR dbg_mem_addr[20] sky130_fd_sc_hd__clkbuf_4
XTAP_6021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput64 net64 VGND VGND VPWR VPWR dbg_mem_addr[30] sky130_fd_sc_hd__buf_2
XFILLER_0_101_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput75 net75 VGND VGND VPWR VPWR dbg_pc[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput86 net86 VGND VGND VPWR VPWR dbg_pc[22] sky130_fd_sc_hd__buf_2
XTAP_6054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput97 net97 VGND VGND VPWR VPWR dbg_pc[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_281_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1622_ _0447_ _0448_ _0451_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__and3_1
XFILLER_0_242_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1553_ _0386_ _0370_ _0371_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_249_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1484_ _1058_ _0319_ _0321_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_120_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_254_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2105_ _0746_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_171_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2036_ _0759_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1076 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer8 net181 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1605_ _0436_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2585_ net142 VGND VGND VPWR VPWR _2585_/X sky130_fd_sc_hd__buf_2
XFILLER_0_239_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1536_ _0336_ _0348_ _0366_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_11_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_279_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1467_ _0954_ _1054_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__nor2_1
XFILLER_0_281_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1398_ _0967_ _0978_ _0996_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_138_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2019_ _0758_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold160 _0214_ VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold171 RF.regs\[1\]\[18\] VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_264_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold182 RF.regs\[1\]\[15\] VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold193 RF.regs\[1\]\[3\] VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1027 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1071 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_267_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2370_ clknet_leaf_4_clk net386 _0168_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1020 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1321_ _0903_ _0934_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__and2b_1
XFILLER_0_276_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1252_ net305 _0897_ _0883_ _0898_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1183_ RF.regs\[1\]\[18\] _0862_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__and2_1
XFILLER_0_190_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2568_ net117 VGND VGND VPWR VPWR _2568_/X sky130_fd_sc_hd__buf_2
XFILLER_0_26_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1519_ ID_EX.ex_rt_data\[9\] net135 net181 VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_273_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2499_ net87 VGND VGND VPWR VPWR _2499_/X sky130_fd_sc_hd__buf_2
XFILLER_0_255_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_266_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1870_ net61 VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__inv_2
XFILLER_0_210_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_255_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2353_ clknet_leaf_15_clk net343 _0151_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_257_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1304_ net79 net78 _0904_ net80 VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__a31o_1
XFILLER_0_252_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2284_ clknet_leaf_11_clk net268 _0082_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1235_ net215 _0895_ _0864_ _0894_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__a22o_1
XFILLER_0_237_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1166_ RF.regs\[1\]\[25\] _0004_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__and2_1
XFILLER_0_189_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1097_ _0823_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1999_ _0756_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_255_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_268_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_261_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1922_ _0634_ _0733_ _0735_ _0585_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__a211o_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1853_ net123 ID_EX.ex_rs_data\[27\] _0591_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1784_ _0588_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__xor2_4
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_269_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2405_ clknet_leaf_1_clk _0302_ VGND VGND VPWR VPWR RF.regs\[1\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_284_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2336_ clknet_leaf_2_clk net23 _0134_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_237_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2267_ clknet_leaf_5_clk net232 _0065_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_256_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1218_ _0846_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_211_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2198_ net358 _0795_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1149_ net35 HAZ.if_id_rt\[0\] _0846_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_941 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold31 RF.regs\[1\]\[2\] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold42 _0236_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold53 ID_EX.ex_rs_data\[23\] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold64 _0229_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold75 ID_EX.ex_rs_data\[8\] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold86 _0231_ VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 ID_EX.ex_rt_data\[7\] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_251_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_6 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_266_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2121_ _0767_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer18 _1020_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
X_2052_ _0761_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer29 _0538_ VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_273_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1905_ _0983_ _0716_ _0717_ _0719_ _0585_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__a311o_1
XFILLER_0_128_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1836_ net122 ID_EX.ex_rs_data\[26\] _0591_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1767_ _0588_ _0589_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1698_ _0520_ _0521_ _0524_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_60_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2319_ clknet_leaf_25_clk net5 _0117_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dfrtp_4
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_259_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput8 net8 VGND VGND VPWR VPWR dbg_alu[15] sky130_fd_sc_hd__clkbuf_4
Xoutput10 net10 VGND VGND VPWR VPWR dbg_alu[17] sky130_fd_sc_hd__clkbuf_4
Xoutput21 net21 VGND VGND VPWR VPWR dbg_alu[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput32 net32 VGND VGND VPWR VPWR dbg_alu[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput43 net43 VGND VGND VPWR VPWR dbg_mem_addr[11] sky130_fd_sc_hd__clkbuf_4
XTAP_6000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput54 net54 VGND VGND VPWR VPWR dbg_mem_addr[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_275_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput65 net65 VGND VGND VPWR VPWR dbg_mem_addr[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_274_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput76 net76 VGND VGND VPWR VPWR dbg_pc[12] sky130_fd_sc_hd__clkbuf_4
Xoutput87 net87 VGND VGND VPWR VPWR dbg_pc[23] sky130_fd_sc_hd__buf_2
XFILLER_0_235_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput98 net98 VGND VGND VPWR VPWR dbg_pc[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_179_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1621_ _0447_ _0448_ _0451_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_112_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1552_ _0370_ _0371_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1483_ _0320_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__buf_6
XFILLER_0_103_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2104_ _0765_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2035_ _0759_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_245_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1819_ _0625_ _0638_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer9 _0610_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_1
XFILLER_0_49_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1604_ _0430_ _0431_ _0434_ _0435_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__a211o_1
XFILLER_0_285_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2584_ net29 VGND VGND VPWR VPWR _2584_/X sky130_fd_sc_hd__buf_2
XFILLER_0_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1535_ _0346_ _0364_ _0365_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_240_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1466_ net132 ID_EX.ex_rs_data\[6\] _1012_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1397_ _0974_ _0977_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__nand2_1
XFILLER_0_207_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2018_ _0758_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold150 ID_EX.ex_rt_data\[26\] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold161 ID_EX.ex_rs_data\[2\] VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold172 RF.regs\[1\]\[10\] VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold183 RF.regs\[1\]\[24\] VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_273_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold194 RF.regs\[1\]\[23\] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1039 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1083 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_249_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1320_ net103 net102 _0902_ net74 VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1251_ net311 _0897_ _0882_ _0898_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__a22o_1
XFILLER_0_276_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_246_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1182_ net245 _0865_ _0870_ _0868_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2567_ net116 VGND VGND VPWR VPWR _2567_/X sky130_fd_sc_hd__buf_2
XFILLER_0_80_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1518_ _1000_ net72 VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2498_ net86 VGND VGND VPWR VPWR _2498_/X sky130_fd_sc_hd__buf_2
XFILLER_0_255_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1449_ _0838_ _1012_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_281_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_270_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_216_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1014 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_269_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2352_ clknet_leaf_15_clk net381 _0150_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1303_ net81 _0905_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__xor2_1
XFILLER_0_270_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2283_ clknet_leaf_11_clk net266 _0081_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_257_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1234_ net292 _0895_ _0863_ _0894_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__a22o_1
XFILLER_0_223_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1165_ net278 _0853_ _0860_ _0855_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_273_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1096_ _0811_ MEM_WB.wb_alu_result\[20\] VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1998_ _0756_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_9011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1921_ _0634_ _0734_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1852_ _0665_ _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_71_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1783_ _0546_ _0602_ _0604_ _0585_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2404_ clknet_leaf_1_clk _0301_ VGND VGND VPWR VPWR RF.regs\[1\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2335_ clknet_leaf_8_clk net22 _0133_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_271_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2266_ clknet_leaf_7_clk net325 _0064_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1217_ net317 _0878_ _0889_ _0881_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__a22o_1
XFILLER_0_237_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2197_ _0748_ net124 _0773_ _0804_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__a31o_1
XFILLER_0_240_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1148_ _0850_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1079_ _0814_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_263_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold32 RF.regs\[1\]\[1\] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold43 ID_EX.ex_rt_data\[20\] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold54 _0268_ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold65 ID_EX.ex_rs_data\[25\] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_243_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold76 _0253_ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold87 ID_EX.ex_rs_data\[14\] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold98 _0220_ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_7 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2120_ _0767_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2051_ _0761_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__inv_2
XFILLER_0_261_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer19 _0955_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_1
XFILLER_0_222_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1904_ _0315_ _0718_ _0634_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1835_ _0640_ _0653_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__xor2_2
XFILLER_0_26_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1766_ _0538_ _0568_ _0587_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1697_ _0315_ _0517_ _0380_ _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__o31a_1
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ clknet_leaf_27_clk net4 _0116_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dfrtp_4
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2249_ clknet_leaf_10_clk net306 _0047_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput11 net11 VGND VGND VPWR VPWR dbg_alu[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_259_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput9 net9 VGND VGND VPWR VPWR dbg_alu[16] sky130_fd_sc_hd__buf_2
Xoutput22 net22 VGND VGND VPWR VPWR dbg_alu[28] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput33 net33 VGND VGND VPWR VPWR dbg_alu[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput44 net44 VGND VGND VPWR VPWR dbg_mem_addr[12] sky130_fd_sc_hd__clkbuf_4
XTAP_6012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput55 net55 VGND VGND VPWR VPWR dbg_mem_addr[22] sky130_fd_sc_hd__clkbuf_4
XTAP_6023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput66 net66 VGND VGND VPWR VPWR dbg_mem_addr[3] sky130_fd_sc_hd__buf_2
XFILLER_0_274_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput77 net77 VGND VGND VPWR VPWR dbg_pc[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput88 net88 VGND VGND VPWR VPWR dbg_pc[24] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_235_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput99 net99 VGND VGND VPWR VPWR dbg_pc[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_200_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_240_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_246_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1620_ _0432_ _0449_ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1551_ _0379_ _0385_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__xor2_2
XFILLER_0_238_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1482_ _1009_ _1040_ _1057_ _0319_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__and4_1
XFILLER_0_254_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_254_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2103_ _0765_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__inv_2
XFILLER_0_222_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2034_ _0759_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1818_ _0634_ _0635_ _0637_ _0585_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1749_ _0432_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_978 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_948 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_250_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_262_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_270_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1603_ _0432_ _0425_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2583_ net28 VGND VGND VPWR VPWR _2583_/X sky130_fd_sc_hd__buf_2
XFILLER_0_10_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1534_ _0369_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1465_ _1058_ _1059_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1396_ _0993_ _0994_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__or2b_1
XFILLER_0_275_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2017_ _0753_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__buf_4
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold140 _0213_ VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold151 _0239_ VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold162 _0247_ VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold173 RF.regs\[1\]\[19\] VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold184 RF.regs\[1\]\[29\] VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_257_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold195 net43 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_273_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_1095 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_243_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1250_ net221 _0897_ _0880_ _0898_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__a22o_1
XFILLER_0_272_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1181_ RF.regs\[1\]\[19\] _0862_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__and2_1
XFILLER_0_215_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2566_ net114 VGND VGND VPWR VPWR _2566_/X sky130_fd_sc_hd__buf_2
XFILLER_0_112_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1517_ _1021_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2497_ net85 VGND VGND VPWR VPWR _2497_/X sky130_fd_sc_hd__buf_2
XFILLER_0_199_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1448_ _1009_ _1025_ _1043_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_177_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1379_ _0967_ net189 ID_EX.ex_aluop\[0\] VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__o21a_1
XFILLER_0_241_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1062 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2351_ clknet_leaf_13_clk net353 _0149_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1302_ _0906_ _0923_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__nor2_1
XFILLER_0_237_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2282_ clknet_leaf_10_clk net316 _0080_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1233_ _0846_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_272_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1164_ RF.regs\[1\]\[26\] _0004_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1095_ _0822_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_4
XFILLER_0_137_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1997_ _0756_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2549_ net126 VGND VGND VPWR VPWR _2549_/X sky130_fd_sc_hd__buf_2
XFILLER_0_239_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_254_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_242_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_249_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_266_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1920_ ID_EX.ex_rt_data\[31\] net128 _0563_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1851_ _0634_ _0666_ _0668_ _0585_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__a211o_2
XFILLER_0_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_976 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_170 VGND VGND VPWR VPWR cpu_top_170/HI dbg_pc[1] sky130_fd_sc_hd__conb_1
XFILLER_0_181_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1782_ _0546_ _0603_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2403_ clknet_leaf_1_clk _0300_ VGND VGND VPWR VPWR RF.regs\[1\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2334_ clknet_leaf_7_clk net21 _0132_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_196_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2265_ clknet_leaf_4_clk net220 _0063_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1216_ RF.regs\[1\]\[3\] _0849_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__and2_1
X_2196_ net362 _0795_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__and2_1
XFILLER_0_237_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1147_ _0844_ net36 _0004_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1078_ _0811_ MEM_WB.wb_alu_result\[29\] VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__and2b_1
XFILLER_0_133_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold33 RF.regs\[1\]\[0\] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_259_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold44 _0233_ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold55 ID_EX.ex_rt_data\[14\] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold66 _0270_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold77 ID_EX.ex_rt_data\[6\] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_243_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold88 _0259_ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold99 ID_EX.ex_rs_data\[21\] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_8 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2050_ _0753_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_221_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1016 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1903_ net64 VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__inv_2
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1834_ _0585_ _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__or2b_1
XFILLER_0_143_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1765_ _0538_ _0568_ _0587_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__or3_4
XFILLER_0_29_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1696_ _0954_ _0522_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__nand2_1
XFILLER_0_269_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2317_ clknet_leaf_9_clk net3 _0115_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dfrtp_4
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ clknet_leaf_10_clk net270 _0046_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_224_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2179_ _0768_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__buf_2
XFILLER_0_240_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput12 net12 VGND VGND VPWR VPWR dbg_alu[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput23 net23 VGND VGND VPWR VPWR dbg_alu[29] sky130_fd_sc_hd__clkbuf_4
Xoutput34 net34 VGND VGND VPWR VPWR dbg_instr[12] sky130_fd_sc_hd__clkbuf_4
Xoutput45 net45 VGND VGND VPWR VPWR dbg_mem_addr[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_274_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput56 net56 VGND VGND VPWR VPWR dbg_mem_addr[23] sky130_fd_sc_hd__buf_2
XFILLER_0_248_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput67 net67 VGND VGND VPWR VPWR dbg_mem_addr[4] sky130_fd_sc_hd__clkbuf_4
XTAP_6035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput78 net78 VGND VGND VPWR VPWR dbg_pc[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput89 net89 VGND VGND VPWR VPWR dbg_pc[25] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_275_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1060 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_240_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1550_ _0380_ _0382_ _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1481_ _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2102_ _0765_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__inv_2
XFILLER_0_253_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2033_ _0759_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1817_ _0546_ _0636_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1748_ _0491_ _0571_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_285_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1679_ _0432_ _0500_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1602_ _0432_ _0433_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_246_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2582_ net27 VGND VGND VPWR VPWR _2582_/X sky130_fd_sc_hd__buf_2
XFILLER_0_281_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1533_ _0352_ _0367_ _0368_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__and3_1
XFILLER_0_267_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1464_ _1009_ _1040_ _1057_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_254_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1395_ _0989_ _0992_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_253_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2016_ _0757_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold130 _0216_ VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold141 ID_EX.ex_rs_data\[10\] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold152 ID_EX.ex_rs_data\[4\] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_257_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold163 ID_EX.ex_rs_data\[5\] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 RF.regs\[1\]\[8\] VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold185 RF.regs\[1\]\[14\] VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold196 net47 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1180_ net253 _0865_ _0869_ _0868_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__a22o_1
XFILLER_0_200_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2565_ net113 VGND VGND VPWR VPWR _2565_/X sky130_fd_sc_hd__buf_2
XFILLER_0_207_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1516_ ID_EX.ex_aluop\[0\] VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2496_ net84 VGND VGND VPWR VPWR _2496_/X sky130_fd_sc_hd__buf_2
XFILLER_0_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1447_ _1042_ _1036_ _1038_ _1039_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__o31a_1
XFILLER_0_215_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1378_ _0974_ _0977_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_156_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_246_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2350_ clknet_leaf_15_clk net383 _0148_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_249_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1301_ net380 _0905_ net82 VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_236_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2281_ clknet_leaf_9_clk net320 _0079_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_237_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1232_ net219 _0890_ _0861_ _0894_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_223_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_1_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_193_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1163_ net257 _0853_ _0859_ _0855_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1094_ _0811_ MEM_WB.wb_alu_result\[21\] VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__and2b_1
XFILLER_0_177_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1996_ _0756_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2548_ net115 VGND VGND VPWR VPWR _2548_/X sky130_fd_sc_hd__buf_2
XFILLER_0_11_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_239_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2479_ net97 VGND VGND VPWR VPWR _2479_/X sky130_fd_sc_hd__buf_2
XFILLER_0_270_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_233_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_231_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_9035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1850_ _0634_ _0667_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_160 VGND VGND VPWR VPWR cpu_top_160/HI dbg_instr[20] sky130_fd_sc_hd__conb_1
XFILLER_0_170_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcpu_top_171 VGND VGND VPWR VPWR cpu_top_171/HI dbg_wb_rd[2] sky130_fd_sc_hd__conb_1
XFILLER_0_280_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1781_ ID_EX.ex_rt_data\[23\] net119 _0563_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_268_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2402_ clknet_leaf_0_clk _0299_ VGND VGND VPWR VPWR RF.regs\[1\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2333_ clknet_leaf_7_clk net20 _0131_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2264_ clknet_leaf_5_clk net293 _0062_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1215_ net326 _0878_ _0888_ _0881_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__a22o_1
XFILLER_0_237_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2195_ _0748_ net123 _0773_ _0803_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1146_ _0849_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1077_ _0813_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_668 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1979_ _0754_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold34 ID.CU.ctrl_alusrc VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold45 ID_EX.ex_rt_data\[25\] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold56 _0227_ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_242_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold67 ID_EX.ex_rt_data\[17\] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold78 _0219_ VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold89 ID_EX.ex_rs_data\[22\] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_9 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_205_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_261_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1028 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1902_ net127 _0563_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1833_ _0383_ net59 _0634_ _0651_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__a31o_1
XFILLER_0_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1764_ _0586_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1695_ net113 ID_EX.ex_rs_data\[18\] _1012_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_271_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ clknet_leaf_12_clk net33 _0114_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dfrtp_4
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2247_ clknet_leaf_10_clk net272 _0045_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_256_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2178_ _0788_ net114 _0786_ _0794_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1129_ _0839_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__inv_4
XFILLER_0_95_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_285_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput13 net13 VGND VGND VPWR VPWR dbg_alu[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput24 net24 VGND VGND VPWR VPWR dbg_alu[2] sky130_fd_sc_hd__clkbuf_4
Xoutput35 net35 VGND VGND VPWR VPWR dbg_instr[16] sky130_fd_sc_hd__buf_2
Xoutput46 net46 VGND VGND VPWR VPWR dbg_mem_addr[14] sky130_fd_sc_hd__clkbuf_4
XTAP_6003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput57 net57 VGND VGND VPWR VPWR dbg_mem_addr[24] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_274_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput68 net68 VGND VGND VPWR VPWR dbg_mem_addr[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_179_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput79 net79 VGND VGND VPWR VPWR dbg_pc[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_200_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_285_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1480_ _1021_ _1070_ _0317_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__o21a_1
XFILLER_0_265_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2101_ _0765_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2032_ _0759_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1816_ ID_EX.ex_rt_data\[25\] net121 _0563_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1747_ net117 ID_EX.ex_rs_data\[21\] _0381_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_269_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1678_ net112 ID_EX.ex_rs_data\[17\] _0381_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_285_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_256_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_263_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_246_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_246_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1601_ net108 ID_EX.ex_rs_data\[13\] _0381_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_242_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2581_ net24 VGND VGND VPWR VPWR _2581_/X sky130_fd_sc_hd__buf_2
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1532_ _0346_ _0349_ _0366_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1463_ _1009_ _1040_ _1057_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1394_ _0989_ _0992_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__and2_1
XFILLER_0_219_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2015_ _0757_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold120 ID_EX.ex_rt_data\[31\] VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 ID_EX.ex_rt_data\[9\] VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold142 _0255_ VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold153 _0249_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold164 RF.regs\[1\]\[30\] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 RF.regs\[1\]\[16\] VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 RF.regs\[1\]\[22\] VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold197 RF.regs\[1\]\[9\] VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_249_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_270_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_259_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2564_ net112 VGND VGND VPWR VPWR _2564_/X sky130_fd_sc_hd__buf_2
XFILLER_0_3_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1515_ _0351_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_254_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2495_ net83 VGND VGND VPWR VPWR _2495_/X sky130_fd_sc_hd__buf_2
XFILLER_0_259_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1446_ _1034_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__buf_4
XFILLER_0_254_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1377_ _0951_ _0975_ _0976_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_278_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1300_ _0907_ _0922_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__nor2_1
XFILLER_0_178_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2280_ clknet_leaf_10_clk net250 _0078_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_252_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1231_ net324 _0890_ _0860_ _0894_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__a22o_1
XFILLER_0_236_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1162_ RF.regs\[1\]\[27\] _0004_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1093_ _0821_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1995_ _0753_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__buf_4
XFILLER_0_117_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2547_ net104 VGND VGND VPWR VPWR _2547_/X sky130_fd_sc_hd__buf_2
XFILLER_0_239_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2478_ net94 VGND VGND VPWR VPWR _2478_/X sky130_fd_sc_hd__buf_2
XFILLER_0_255_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_270_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1429_ net202 net186 VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_208_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcpu_top_150 VGND VGND VPWR VPWR cpu_top_150/HI dbg_instr[8] sky130_fd_sc_hd__conb_1
XFILLER_0_86_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcpu_top_161 VGND VGND VPWR VPWR cpu_top_161/HI dbg_instr[22] sky130_fd_sc_hd__conb_1
XFILLER_0_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1780_ _0383_ net56 VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_172 VGND VGND VPWR VPWR cpu_top_172/HI dbg_wb_rd[3] sky130_fd_sc_hd__conb_1
XFILLER_0_170_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2401_ clknet_leaf_1_clk _0298_ VGND VGND VPWR VPWR RF.regs\[1\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2332_ clknet_leaf_8_clk net139 _0130_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2263_ clknet_leaf_3_clk net216 _0061_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1214_ RF.regs\[1\]\[4\] _0849_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2194_ net354 _0795_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__and2_1
XFILLER_0_215_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1145_ _0846_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__inv_2
XFILLER_0_250_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1076_ _0811_ MEM_WB.wb_alu_result\[30\] VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1978_ _0754_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold35 RF.regs\[1\]\[4\] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold46 _0238_ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold57 ID_EX.ex_rt_data\[27\] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold68 _0230_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold79 ID_EX.ex_rs_data\[20\] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_978 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1901_ ID_EX.ex_rt_data\[30\] net199 VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1832_ ID_EX.ex_rt_data\[26\] _0563_ _0650_ _0983_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1763_ _0546_ _0582_ _0584_ _0585_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_269_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1694_ _0403_ _0466_ _0504_ _0519_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_40_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2315_ clknet_leaf_13_clk net32 _0113_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfrtp_4
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ clknet_leaf_10_clk net252 _0044_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_224_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2177_ net347 _0782_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1128_ MEM_WB.wb_memtoreg MEM_WB.wb_alu_result\[4\] VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__or2b_2
XFILLER_0_79_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_285_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput14 net140 VGND VGND VPWR VPWR dbg_alu[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_202_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput25 net25 VGND VGND VPWR VPWR dbg_alu[30] sky130_fd_sc_hd__buf_4
XFILLER_0_47_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput36 net36 VGND VGND VPWR VPWR dbg_instr[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput47 net47 VGND VGND VPWR VPWR dbg_mem_addr[15] sky130_fd_sc_hd__clkbuf_4
XTAP_6015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput58 net58 VGND VGND VPWR VPWR dbg_mem_addr[25] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput69 net69 VGND VGND VPWR VPWR dbg_mem_addr[6] sky130_fd_sc_hd__buf_2
XFILLER_0_124_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_281_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2100_ _0765_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2031_ _0759_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__inv_2
XFILLER_0_206_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1815_ _0383_ net58 VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_245_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1746_ _0538_ _0550_ _0567_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1677_ _0488_ _0503_ _0504_ _0473_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_284_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2229_ clknet_leaf_19_clk _0203_ _0027_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_280_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1600_ _1011_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__clkbuf_4
X_2580_ net13 VGND VGND VPWR VPWR _2580_/X sky130_fd_sc_hd__buf_2
XFILLER_0_124_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1531_ _0346_ _0349_ _0366_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__or3_1
XFILLER_0_267_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1462_ _1056_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1393_ _0951_ _0986_ _0991_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_250_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2014_ _0757_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold110 ID_EX.ex_rt_data\[13\] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _0244_ VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1729_ _0432_ _0552_ _0553_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__o21ai_1
Xhold132 _0222_ VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold143 ID_EX.ex_rs_data\[3\] VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 ID_EX.ex_rt_data\[4\] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold165 ID_EX.ex_rt_data\[2\] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold176 RF.regs\[1\]\[11\] VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold187 RF.regs\[1\]\[25\] VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold198 net72 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2563_ net111 VGND VGND VPWR VPWR _2563_/X sky130_fd_sc_hd__buf_2
XFILLER_0_207_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1514_ _0349_ ID_EX.ex_aluop\[0\] _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__and3b_1
XFILLER_0_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2494_ net82 VGND VGND VPWR VPWR _2494_/X sky130_fd_sc_hd__buf_2
XFILLER_0_107_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1445_ _1009_ _1040_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1376_ _0951_ _0971_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_235_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_249_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1230_ net231 _0890_ _0859_ _0894_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1161_ net286 _0853_ _0858_ _0855_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__a22o_1
XFILLER_0_251_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_254_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1092_ _0810_ MEM_WB.wb_alu_result\[22\] VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__and2b_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_250_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1994_ _0755_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2615_ net73 VGND VGND VPWR VPWR _2615_/X sky130_fd_sc_hd__buf_2
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2546_ net65 VGND VGND VPWR VPWR _2546_/X sky130_fd_sc_hd__buf_2
XFILLER_0_122_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1428_ _1021_ _1022_ _1024_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_254_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1359_ net137 net138 FU.id_ex_rt\[0\] net136 VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__and4b_2
XFILLER_0_39_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire139 net19 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_4
XFILLER_0_135_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_151 VGND VGND VPWR VPWR cpu_top_151/HI dbg_instr[9] sky130_fd_sc_hd__conb_1
XFILLER_0_167_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_162 VGND VGND VPWR VPWR cpu_top_162/HI dbg_instr[23] sky130_fd_sc_hd__conb_1
XFILLER_0_0_1631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_173 VGND VGND VPWR VPWR cpu_top_173/HI dbg_wb_rd[4] sky130_fd_sc_hd__conb_1
XFILLER_0_154_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2400_ clknet_leaf_5_clk _0297_ VGND VGND VPWR VPWR RF.regs\[1\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_268_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2331_ clknet_leaf_4_clk net18 _0129_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_62_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2262_ clknet_leaf_5_clk net234 _0060_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_236_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1213_ net337 _0878_ _0887_ _0881_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2193_ _0748_ net122 _0773_ _0802_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1144_ _0848_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_251_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1075_ _0812_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_250_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1977_ _0754_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2529_ net46 VGND VGND VPWR VPWR _2529_/X sky130_fd_sc_hd__buf_2
XFILLER_0_80_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold36 RF.regs\[1\]\[5\] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold47 ID_EX.ex_rt_data\[11\] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_270_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold58 _0240_ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold69 ID_EX.ex_rs_data\[24\] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_268_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1900_ _0715_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_4
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1831_ net122 net199 VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1762_ _1042_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1693_ _0403_ _0466_ _0504_ _0519_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2314_ clknet_leaf_14_clk net31 _0112_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dfrtp_4
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2245_ clknet_leaf_9_clk _0218_ _0043_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_206_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2176_ _0788_ net113 _0786_ _0793_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1127_ _0838_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__inv_2
XFILLER_0_221_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput15 net15 VGND VGND VPWR VPWR dbg_alu[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_247_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput26 net26 VGND VGND VPWR VPWR dbg_alu[31] sky130_fd_sc_hd__buf_8
XFILLER_0_222_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput37 net37 VGND VGND VPWR VPWR dbg_instr[26] sky130_fd_sc_hd__clkbuf_4
XTAP_6005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput48 net48 VGND VGND VPWR VPWR dbg_mem_addr[16] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_247_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput59 net59 VGND VGND VPWR VPWR dbg_mem_addr[26] sky130_fd_sc_hd__buf_2
XTAP_6016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_268_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_285_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_266_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2030_ _0759_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__inv_2
XTAP_5893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1814_ _0546_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__buf_2
XFILLER_0_2_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1745_ net333 _0568_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_269_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1676_ _0487_ _0503_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_245_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2228_ clknet_leaf_19_clk _0202_ _0026_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_240_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2159_ net350 _0782_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__and2_1
XFILLER_0_240_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1530_ _0364_ _0365_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1461_ _1021_ _1053_ _1055_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__o21a_1
XFILLER_0_227_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1392_ _0841_ net193 _0990_ _0954_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__o211a_1
XFILLER_0_279_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_253_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2013_ _0757_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__inv_2
XFILLER_0_261_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold100 _0266_ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold111 _0226_ VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1728_ _0432_ _0548_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__nand2_1
Xhold122 ID_EX.ex_rs_data\[7\] VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold133 ID_EX.ex_rs_data\[30\] VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold144 _0248_ VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold155 _0217_ VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _0215_ VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold177 RF.regs\[1\]\[20\] VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ _0403_ _0466_ _0487_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold188 RF.regs\[1\]\[28\] VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold199 net54 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_896 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2562_ net110 VGND VGND VPWR VPWR _2562_/X sky130_fd_sc_hd__buf_2
XFILLER_0_140_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1513_ _0336_ _0348_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2493_ net81 VGND VGND VPWR VPWR _2493_/X sky130_fd_sc_hd__buf_2
XFILLER_0_103_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_16
X_1444_ _1034_ _1036_ _1038_ _1025_ _1039_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__o311a_4
XFILLER_0_43_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1375_ net115 ID_EX.ex_rs_data\[1\] _0955_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_253_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_242_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_246_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_671 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_249_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1160_ RF.regs\[1\]\[28\] _0004_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__and2_1
XFILLER_0_159_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1091_ _0820_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_4
XTAP_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1993_ _0755_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2614_ net39 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
XFILLER_0_70_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2545_ net64 VGND VGND VPWR VPWR _2545_/X sky130_fd_sc_hd__buf_2
XFILLER_0_267_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1427_ _1021_ _1023_ EX_MEM.ex_memread VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_177_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1358_ _0958_ _0951_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__nand2_1
XFILLER_0_272_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1289_ net89 _0910_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_285_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_152 VGND VGND VPWR VPWR cpu_top_152/HI dbg_instr[10] sky130_fd_sc_hd__conb_1
XFILLER_0_0_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_249_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcpu_top_163 VGND VGND VPWR VPWR cpu_top_163/HI dbg_instr[24] sky130_fd_sc_hd__conb_1
XFILLER_0_37_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_674 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2330_ clknet_leaf_3_clk net17 _0128_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2261_ clknet_leaf_2_clk net226 _0059_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1212_ RF.regs\[1\]\[5\] _0875_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__and2_1
XFILLER_0_251_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2192_ net355 _0795_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1143_ net39 ID.CU.ctrl_alusrc _0846_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1074_ _0811_ MEM_WB.wb_alu_result\[31\] VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__and2b_1
XFILLER_0_220_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1976_ _0754_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_268_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2528_ net45 VGND VGND VPWR VPWR _2528_/X sky130_fd_sc_hd__buf_2
XFILLER_0_122_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold37 _0286_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold48 _0224_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold59 ID_EX.ex_rt_data\[22\] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_8178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1830_ _0647_ _0648_ _0649_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1761_ _0546_ _0583_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1692_ _0983_ _0515_ _0516_ _0518_ _1042_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__a311o_1
XFILLER_0_282_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2313_ clknet_leaf_9_clk net30 _0111_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dfrtp_4
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2244_ clknet_leaf_16_clk net329 _0042_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_206_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2175_ net345 _0782_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1126_ _0809_ MEM_WB.wb_alu_result\[5\] VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_36_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1959_ _0751_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput16 net16 VGND VGND VPWR VPWR dbg_alu[22] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_275_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput27 net27 VGND VGND VPWR VPWR dbg_alu[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput38 net38 VGND VGND VPWR VPWR dbg_instr[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput49 net49 VGND VGND VPWR VPWR dbg_mem_addr[17] sky130_fd_sc_hd__clkbuf_4
XTAP_6006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_285_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_285_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_251_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1813_ _0620_ _0632_ _0633_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__o21a_2
XFILLER_0_155_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1744_ _0550_ _0567_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1675_ _0390_ _0500_ _0502_ _1042_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__a211o_1
XFILLER_0_284_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2227_ clknet_leaf_19_clk _0201_ _0025_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_213_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2158_ _0005_ net105 _0774_ _0783_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1109_ _0829_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_6
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2089_ _0764_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__inv_2
XFILLER_0_269_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_276_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1028 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1460_ _1021_ _1054_ EX_MEM.ex_memread VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_266_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_266_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1391_ ID_EX.ex_rs_data\[2\] net193 VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__nand2_1
XFILLER_0_285_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_282_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2012_ _0757_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold101 ID_EX.ex_rs_data\[0\] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold112 ID_EX.ex_rs_data\[28\] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1727_ net116 ID_EX.ex_rs_data\[20\] _0381_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold123 _0252_ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold134 _0275_ VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold145 ID_EX.ex_rs_data\[9\] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold156 ID_EX.ex_rt_data\[30\] VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_284_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold167 RF.regs\[1\]\[12\] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ _0390_ _0484_ _0486_ _1034_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__a211o_1
XFILLER_0_258_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold178 RF.regs\[1\]\[17\] VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_284_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold189 RF.regs\[1\]\[31\] VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1589_ _0413_ _0421_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__nor2_1
XFILLER_0_238_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_241_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2561_ net109 VGND VGND VPWR VPWR _2561_/X sky130_fd_sc_hd__buf_2
XFILLER_0_144_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1512_ _0336_ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2492_ net80 VGND VGND VPWR VPWR _2492_/X sky130_fd_sc_hd__buf_2
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1443_ ID_EX.ex_imm\[12\] _1034_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_227_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_259_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1374_ _0966_ _0973_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_235_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1027 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1090_ _0811_ MEM_WB.wb_alu_result\[23\] VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__and2b_1
XFILLER_0_137_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1992_ _0755_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2613_ net39 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_259_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2544_ net62 VGND VGND VPWR VPWR _2544_/X sky130_fd_sc_hd__buf_2
XFILLER_0_140_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1426_ net73 net67 VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__or2b_1
XFILLER_0_254_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1357_ net73 net41 VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__nor2_1
XFILLER_0_270_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1288_ net384 _0911_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_153 VGND VGND VPWR VPWR cpu_top_153/HI dbg_instr[11] sky130_fd_sc_hd__conb_1
Xcpu_top_164 VGND VGND VPWR VPWR cpu_top_164/HI dbg_instr[25] sky130_fd_sc_hd__conb_1
XFILLER_0_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_283_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2260_ clknet_leaf_2_clk net218 _0058_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_236_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1211_ net282 _0878_ _0886_ _0881_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_284_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2191_ _0748_ net121 _0773_ _0801_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1142_ _0847_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1073_ _0810_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_254_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1975_ _0754_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2527_ net44 VGND VGND VPWR VPWR _2527_/X sky130_fd_sc_hd__buf_2
XFILLER_0_268_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold38 EX_MEM.mem_regwrite VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ _0982_ _0985_ _0987_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__a21o_1
XFILLER_0_215_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold49 ID_EX.ex_rt_data\[15\] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ clknet_leaf_9_clk net211 VGND VGND VPWR VPWR RF.regs\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1760_ ID_EX.ex_rt_data\[22\] net118 _0373_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1691_ _0315_ _0517_ _0390_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_204_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2312_ clknet_leaf_14_clk net29 _0110_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dfrtp_4
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2243_ clknet_leaf_16_clk net304 _0041_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2174_ _0788_ net112 _0786_ _0792_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__a31o_1
XFILLER_0_215_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1125_ _0837_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_221_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1958_ _0751_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__inv_2
XFILLER_0_181_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1889_ _0684_ _0689_ _0703_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput17 net17 VGND VGND VPWR VPWR dbg_alu[23] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput28 net28 VGND VGND VPWR VPWR dbg_alu[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_222_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput39 net39 VGND VGND VPWR VPWR dbg_instr[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_247_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1812_ _0620_ _0632_ _0980_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1743_ _0546_ _0564_ _0566_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1674_ _0353_ _0501_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2226_ clknet_leaf_19_clk _0200_ _0024_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_253_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2157_ net346 _0782_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__and2_1
XFILLER_0_273_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1108_ _0810_ MEM_WB.wb_alu_result\[14\] VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2088_ _0764_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1035 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_278_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1390_ _0981_ _0988_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_281_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_250_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2011_ _0757_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1726_ net333 _0550_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__xnor2_2
Xhold102 ID_EX.ex_rs_data\[29\] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold113 _0273_ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_258_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold124 ID_EX.ex_rt_data\[28\] VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold135 ID_EX.ex_rs_data\[15\] VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold146 _0254_ VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__dlygate4sd3_1
X_1657_ _0353_ _0485_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold157 _0243_ VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_285_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold168 RF.regs\[1\]\[13\] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 net68 VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1588_ _0417_ _0420_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2209_ clknet_leaf_15_clk _0183_ _0007_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_252_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2560_ net108 VGND VGND VPWR VPWR _2560_/X sky130_fd_sc_hd__buf_2
XFILLER_0_84_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1511_ _0346_ _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2491_ net79 VGND VGND VPWR VPWR _2491_/X sky130_fd_sc_hd__buf_2
XFILLER_0_80_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1442_ _1021_ _1037_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__and2_1
XFILLER_0_266_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1373_ _0964_ _0970_ _0972_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_219_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_270_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_832 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1039 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1709_ _0390_ _0534_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__nor2_1
XFILLER_0_258_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1991_ _0755_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2612_ net36 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_246_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2543_ net61 VGND VGND VPWR VPWR _2543_/X sky130_fd_sc_hd__buf_2
XFILLER_0_100_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1425_ ID_EX.ex_rt_data\[4\] net130 _1003_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__mux2_4
XFILLER_0_259_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1356_ _0951_ _0956_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__or2_1
XFILLER_0_253_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1287_ _0912_ _0917_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_231_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_285_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_143 VGND VGND VPWR VPWR cpu_top_143/HI dbg_instr[0] sky130_fd_sc_hd__conb_1
XFILLER_0_182_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcpu_top_154 VGND VGND VPWR VPWR cpu_top_154/HI dbg_instr[13] sky130_fd_sc_hd__conb_1
XFILLER_0_65_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcpu_top_165 VGND VGND VPWR VPWR cpu_top_165/HI dbg_instr[28] sky130_fd_sc_hd__conb_1
XFILLER_0_282_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_268_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1210_ RF.regs\[1\]\[6\] _0875_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2190_ net361 _0795_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__and2_1
XFILLER_0_178_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1141_ _0844_ FU.id_ex_rs\[0\] _0846_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_260_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1072_ _0809_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1974_ _0754_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2526_ net43 VGND VGND VPWR VPWR _2526_/X sky130_fd_sc_hd__buf_2
XFILLER_0_140_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1408_ _0981_ _0988_ _1005_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__o21ba_1
Xhold39 net71 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_270_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2388_ clknet_leaf_16_clk _0285_ VGND VGND VPWR VPWR RF.regs\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1339_ _0900_ _0945_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_838 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1690_ net50 VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_243_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2311_ clknet_leaf_14_clk net28 _0109_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dfrtp_4
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2242_ clknet_leaf_16_clk net340 _0040_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2173_ net352 _0782_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__and2_1
XFILLER_0_252_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1124_ _0809_ MEM_WB.wb_alu_result\[6\] VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__and2b_1
XFILLER_0_233_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1957_ _0751_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1888_ _0684_ _0689_ _0703_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput18 net18 VGND VGND VPWR VPWR dbg_alu[24] sky130_fd_sc_hd__buf_2
XFILLER_0_275_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput29 net29 VGND VGND VPWR VPWR dbg_alu[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2509_ net36 VGND VGND VPWR VPWR _2509_/X sky130_fd_sc_hd__buf_2
XFILLER_0_25_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_243_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_268_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_249_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_27_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_203_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1811_ _0630_ _0631_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1742_ _0546_ _0565_ _1042_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1673_ ID_EX.ex_rt_data\[17\] net112 _0373_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ clknet_leaf_19_clk _0199_ _0023_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_213_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2156_ _0768_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__buf_2
XFILLER_0_55_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1107_ _0828_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_221_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2087_ _0764_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_18_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2010_ _0757_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1725_ _0546_ _0547_ _0549_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold103 _0274_ VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_285_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold114 ID_EX.ex_rs_data\[18\] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 ID_EX.ex_rs_data\[13\] VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_7_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_16
Xhold136 _0260_ VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1081 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold147 ID_EX.ex_rs_data\[1\] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__dlygate4sd3_1
X_1656_ ID_EX.ex_rt_data\[16\] net111 net181 VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__mux2_1
Xhold158 net50 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_257_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold169 net70 VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_284_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_229_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1587_ _0386_ _0370_ _0399_ _0418_ _0419_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__a311o_1
XFILLER_0_284_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2208_ clknet_leaf_18_clk _0182_ _0006_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2139_ net205 _0769_ _0772_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1510_ _0341_ _0345_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2490_ net78 VGND VGND VPWR VPWR _2490_/X sky130_fd_sc_hd__buf_2
XFILLER_0_224_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1441_ _1000_ net68 VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_259_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1372_ _0964_ _0971_ EX_MEM.ex_memread VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1708_ ID_EX.ex_rt_data\[19\] net114 _0373_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1639_ net110 ID_EX.ex_rs_data\[15\] _1012_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_258_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1990_ _0755_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2611_ net36 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2542_ net60 VGND VGND VPWR VPWR _2542_/X sky130_fd_sc_hd__buf_2
XFILLER_0_49_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1424_ _0964_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__buf_2
XFILLER_0_282_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1355_ net104 ID_EX.ex_rs_data\[0\] _0955_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1286_ net90 _0911_ net91 VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_194_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_270_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_277_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_285_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_277_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_144 VGND VGND VPWR VPWR cpu_top_144/HI dbg_instr[1] sky130_fd_sc_hd__conb_1
Xcpu_top_155 VGND VGND VPWR VPWR cpu_top_155/HI dbg_instr[14] sky130_fd_sc_hd__conb_1
XFILLER_0_182_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_166 VGND VGND VPWR VPWR cpu_top_166/HI dbg_instr[29] sky130_fd_sc_hd__conb_1
XFILLER_0_65_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1668 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1140_ _0845_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_191_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1071_ MEM_WB.wb_memtoreg VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_232_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_267_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1973_ _0753_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__buf_4
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2525_ net42 VGND VGND VPWR VPWR _2525_/X sky130_fd_sc_hd__buf_2
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1407_ _0964_ _1001_ _1002_ _1004_ EX_MEM.ex_memread VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__a221o_1
Xhold29 EX_MEM.ex_regwrite VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_243_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2387_ clknet_leaf_9_clk _0284_ VGND VGND VPWR VPWR RF.regs\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_255_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1338_ net94 _0004_ net97 VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1269_ net77 net76 net75 _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__and4_2
XFILLER_0_272_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2310_ clknet_leaf_15_clk net27 _0108_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dfrtp_4
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2241_ clknet_leaf_16_clk net334 _0039_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_218_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2172_ _0788_ net111 _0786_ _0791_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__a31o_1
XFILLER_0_178_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1123_ _0836_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__buf_4
XFILLER_0_117_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1956_ _0751_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1887_ _0634_ _0700_ _0702_ _0585_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput19 net139 VGND VGND VPWR VPWR dbg_alu[25] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2508_ net36 VGND VGND VPWR VPWR _2508_/X sky130_fd_sc_hd__buf_2
XFILLER_0_274_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_214_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1810_ _0626_ _0629_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1741_ _0343_ net54 VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1672_ _0343_ net49 VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_256_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ clknet_leaf_19_clk _0198_ _0022_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_280_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2155_ _0005_ net135 _0774_ _0781_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1106_ _0810_ MEM_WB.wb_alu_result\[15\] VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2086_ _0764_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1939_ _0749_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__buf_4
XFILLER_0_280_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_250_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1724_ _0390_ _0548_ _1042_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold104 ID_EX.ex_rs_data\[26\] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold115 _0263_ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold126 _0258_ VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1655_ _1000_ net48 VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_258_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold137 ID_EX.ex_rt_data\[10\] VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold148 _0246_ VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1586_ _0395_ _0398_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_258_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2207_ clknet_leaf_8_clk _0181_ _0005_ VGND VGND VPWR VPWR FU.id_ex_rt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_20_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2138_ _0747_ net126 _0953_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2069_ _0762_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__inv_2
XFILLER_0_234_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1008 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_246_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_254_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1440_ _0838_ net196 _1035_ _0982_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__o211a_1
XFILLER_0_266_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1371_ net73 net52 VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__nor2_1
XFILLER_0_282_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_231_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1707_ _0343_ net51 VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__nand2_1
XFILLER_0_281_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1638_ _0402_ _0429_ _0446_ _0464_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1569_ _0321_ _0358_ _0376_ _0394_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__and4_4
XFILLER_0_226_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_257_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2610_ net26 VGND VGND VPWR VPWR _2610_/X sky130_fd_sc_hd__buf_2
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2541_ net59 VGND VGND VPWR VPWR _2541_/X sky130_fd_sc_hd__buf_2
XFILLER_0_183_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_282_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1423_ _0999_ _1017_ _1016_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__a21o_1
XFILLER_0_227_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1354_ FU.id_ex_rs\[0\] _0953_ _0954_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__nand3_4
XFILLER_0_235_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1285_ _0913_ _0916_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__nor2_1
XFILLER_0_250_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_249_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_145 VGND VGND VPWR VPWR cpu_top_145/HI dbg_instr[2] sky130_fd_sc_hd__conb_1
XFILLER_0_64_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_156 VGND VGND VPWR VPWR cpu_top_156/HI dbg_instr[15] sky130_fd_sc_hd__conb_1
XFILLER_0_163_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcpu_top_167 VGND VGND VPWR VPWR cpu_top_167/HI dbg_instr[30] sky130_fd_sc_hd__conb_1
XFILLER_0_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1972_ _0746_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2524_ net72 VGND VGND VPWR VPWR _2524_/X sky130_fd_sc_hd__buf_2
XFILLER_0_60_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1406_ net129 _1003_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__nand2_1
X_2386_ clknet_leaf_16_clk _0283_ VGND VGND VPWR VPWR RF.regs\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_282_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1337_ _0901_ _0944_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__nor2_1
XFILLER_0_236_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1268_ net74 net103 net102 _0902_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__and4_1
XFILLER_0_250_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1199_ RF.regs\[1\]\[11\] _0875_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_277_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ clknet_leaf_16_clk net314 _0038_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2171_ net349 _0782_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1122_ _0809_ MEM_WB.wb_alu_result\[7\] VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__and2b_1
XFILLER_0_156_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1955_ _0751_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1886_ _0634_ _0701_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2507_ net96 VGND VGND VPWR VPWR _2507_/X sky130_fd_sc_hd__buf_2
XFILLER_0_60_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_282_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2369_ clknet_leaf_4_clk net396 _0167_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_285_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_249_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1740_ ID_EX.ex_rt_data\[21\] net117 _0563_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1671_ _0497_ _0483_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__and2b_1
XFILLER_0_159_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2223_ clknet_1_0__leaf_clk _0197_ _0021_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_178_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2154_ net371 _0769_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1105_ _0827_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_6
XFILLER_0_108_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2085_ _0764_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__inv_2
XFILLER_0_220_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1938_ _0746_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1869_ net124 _0563_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1723_ _0343_ net53 VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold105 _0271_ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold116 ID_EX.ex_rt_data\[19\] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold127 ID_EX.ex_rs_data\[31\] VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1654_ _0417_ _0479_ _0480_ _0482_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__a211o_4
XFILLER_0_83_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_262_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold138 _0223_ VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold149 ID_EX.ex_rt_data\[5\] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_273_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1585_ _0395_ _0398_ _0379_ _0385_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_281_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2206_ net97 net94 VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2137_ net206 _0769_ _0771_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__a21o_1
XFILLER_0_221_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2068_ _0762_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__inv_2
XFILLER_0_230_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_246_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1370_ ID_EX.ex_rt_data\[1\] net115 _0960_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__mux2_4
XFILLER_0_281_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_229_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1706_ _0532_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_4
XFILLER_0_170_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1637_ _0403_ _0466_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_258_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1568_ _0399_ _0400_ _0401_ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__a21oi_4
XFILLER_0_26_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1499_ _1068_ _0331_ _0335_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_193_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2540_ net58 VGND VGND VPWR VPWR _2540_/X sky130_fd_sc_hd__buf_2
XFILLER_0_144_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1422_ _0980_ _1019_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__nor2_8
XFILLER_0_239_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_259_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1353_ EX_MEM.mem_rd\[1\] EX_MEM.mem_regwrite FU.id_ex_rs\[0\] EX_MEM.mem_rd\[0\]
+ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_282_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1284_ net92 _0912_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__nor2_1
XFILLER_0_251_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_146 VGND VGND VPWR VPWR cpu_top_146/HI dbg_instr[3] sky130_fd_sc_hd__conb_1
XFILLER_0_110_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_157 VGND VGND VPWR VPWR cpu_top_157/HI dbg_instr[17] sky130_fd_sc_hd__conb_1
XFILLER_0_64_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_168 VGND VGND VPWR VPWR cpu_top_168/HI dbg_memwrite sky130_fd_sc_hd__conb_1
XFILLER_0_184_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_232_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1971_ _0752_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__inv_2
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2523_ net71 VGND VGND VPWR VPWR _2523_/X sky130_fd_sc_hd__buf_2
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1405_ _0960_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__buf_6
XFILLER_0_227_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2385_ clknet_leaf_9_clk _0282_ VGND VGND VPWR VPWR RF.regs\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_283_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1336_ net98 _0900_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_235_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 rst VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
XFILLER_0_251_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1267_ net101 net100 net99 _0901_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__and4_1
XFILLER_0_170_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1198_ net267 _0878_ _0879_ _0868_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_282_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2170_ _0788_ net110 _0786_ _0790_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__a31o_1
XFILLER_0_228_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1121_ _0835_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_233_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1954_ _0751_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1885_ ID_EX.ex_rt_data\[29\] net125 _0563_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2506_ net95 VGND VGND VPWR VPWR _2506_/X sky130_fd_sc_hd__buf_2
XFILLER_0_25_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2368_ clknet_leaf_27_clk net55 _0166_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1319_ _0933_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__clkbuf_1
XTAP_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2299_ clknet_leaf_7_clk net258 _0097_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_251_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_240_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_249_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1670_ _0980_ _0498_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__nor2_4
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ clknet_1_0__leaf_clk _0196_ _0020_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_139_1014 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2153_ _0005_ net134 _0774_ _0780_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__a31o_1
XFILLER_0_108_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1104_ _0809_ MEM_WB.wb_alu_result\[16\] VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__and2b_1
XFILLER_0_152_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2084_ _0764_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_863 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1937_ _0748_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1868_ ID_EX.ex_rt_data\[28\] net199 VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1799_ _0483_ _0557_ _0614_ _0618_ _0619_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__a311o_4
XFILLER_0_275_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_278_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_914 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_268_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1722_ ID_EX.ex_rt_data\[20\] net116 _0373_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold106 ID_EX.ex_rs_data\[16\] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 _0232_ VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1653_ _0454_ _0456_ _0475_ _0481_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__a31o_1
XFILLER_0_13_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold128 _0276_ VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold139 ID_EX.ex_rt_data\[0\] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_262_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1584_ _0414_ _0415_ _0335_ _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__o31a_1
XFILLER_0_201_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_265_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_275_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2205_ _0808_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2136_ _0747_ net115 _0953_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__and3_1
XFILLER_0_178_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2067_ _0762_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_275_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_270_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1705_ _0352_ _0530_ _0531_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1636_ _0465_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__buf_2
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1567_ _0399_ _0400_ _0969_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_285_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1498_ _0327_ _0333_ _0334_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2119_ _0767_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_254_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1421_ net200 _1018_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__xor2_4
XFILLER_0_121_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1352_ _0952_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__buf_2
XFILLER_0_208_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1283_ net93 _0913_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__xor2_1
XFILLER_0_250_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_696 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1619_ _0432_ _0443_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__nand2_1
XTAP_6919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2599_ net140 VGND VGND VPWR VPWR _2599_/X sky130_fd_sc_hd__buf_2
XFILLER_0_26_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcpu_top_147 VGND VGND VPWR VPWR cpu_top_147/HI dbg_instr[4] sky130_fd_sc_hd__conb_1
Xcpu_top_158 VGND VGND VPWR VPWR cpu_top_158/HI dbg_instr[18] sky130_fd_sc_hd__conb_1
XFILLER_0_181_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_169 VGND VGND VPWR VPWR cpu_top_169/HI dbg_pc[0] sky130_fd_sc_hd__conb_1
XFILLER_0_247_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1970_ _0752_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__inv_2
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2522_ net70 VGND VGND VPWR VPWR _2522_/X sky130_fd_sc_hd__buf_2
XFILLER_0_12_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1404_ ID_EX.ex_rt_data\[3\] _0962_ _0964_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2384_ clknet_leaf_16_clk _0281_ VGND VGND VPWR VPWR RF.regs\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1335_ _0943_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_282_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1266_ net98 _0900_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__and2_1
XFILLER_0_237_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1197_ RF.regs\[1\]\[12\] _0875_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_285_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1020 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1120_ _0809_ MEM_WB.wb_alu_result\[8\] VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_267_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_695 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1953_ _0751_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1884_ _0383_ net62 VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2505_ net93 VGND VGND VPWR VPWR _2505_/X sky130_fd_sc_hd__buf_2
XFILLER_0_45_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2367_ clknet_leaf_2_clk net373 _0165_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_236_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1318_ _0931_ _0932_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2298_ clknet_leaf_7_clk net279 _0096_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_212_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1249_ HAZ.if_id_rt\[0\] VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_212_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_220_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_249_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ clknet_leaf_24_clk _0195_ _0019_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_280_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1026 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2152_ net348 _0769_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__and2_1
XFILLER_0_238_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1103_ _0826_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_4
XFILLER_0_108_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2083_ _0746_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__buf_4
XFILLER_0_117_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_271_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1936_ _0747_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_956 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1867_ _0665_ _0669_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__and2_4
XFILLER_0_44_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1798_ _0560_ _0559_ _0595_ _0597_ _0610_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_124_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_278_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_240_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1721_ _0390_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1652_ _0452_ _0474_ _0472_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__a21o_1
Xhold107 _0261_ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold118 ID_EX.ex_rt_data\[24\] VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold129 ID_EX.ex_rt_data\[3\] VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1583_ _0348_ _0366_ _0386_ _0399_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__and4b_1
XFILLER_0_61_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2204_ _0000_ net94 VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__and2_1
XFILLER_0_281_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2135_ net207 _0769_ _0770_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__a21o_1
XFILLER_0_252_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2066_ _0762_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1919_ _0383_ net65 VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_229_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1704_ _0528_ _0529_ _0527_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1635_ _0429_ _0446_ _0464_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__and3_1
XFILLER_0_258_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1566_ _0379_ _0385_ _0387_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1497_ _0322_ _0325_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__or2b_1
XFILLER_0_265_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2118_ _0767_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2049_ _0760_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_265_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1000 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1420_ _1016_ _1017_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__or2b_2
XFILLER_0_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1351_ net137 net177 net136 VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__and3b_1
XFILLER_0_248_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1282_ _0914_ _0915_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__nor2_1
XFILLER_0_263_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_231_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1618_ net109 ID_EX.ex_rs_data\[14\] _0381_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2598_ net12 VGND VGND VPWR VPWR _2598_/X sky130_fd_sc_hd__buf_2
XFILLER_0_22_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1549_ _0383_ net42 _1011_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcpu_top_148 VGND VGND VPWR VPWR cpu_top_148/HI dbg_instr[6] sky130_fd_sc_hd__conb_1
Xcpu_top_159 VGND VGND VPWR VPWR cpu_top_159/HI dbg_instr[19] sky130_fd_sc_hd__conb_1
XFILLER_0_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_268_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2521_ net69 VGND VGND VPWR VPWR _2521_/X sky130_fd_sc_hd__buf_2
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_279_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1403_ _1000_ net66 VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__nand2_1
XFILLER_0_209_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2383_ clknet_leaf_18_clk _0000_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_20_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1334_ _0941_ _0942_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__and2_1
XFILLER_0_237_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1265_ net97 net94 _0849_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__and3_1
XFILLER_0_250_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1196_ _0846_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_231_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1952_ _0751_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__inv_2
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1883_ _0699_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2504_ net92 VGND VGND VPWR VPWR _2504_/X sky130_fd_sc_hd__buf_2
XFILLER_0_109_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_259_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2366_ clknet_leaf_26_clk net399 _0164_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1317_ net75 _0903_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__or2_1
XFILLER_0_224_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2297_ clknet_leaf_4_clk net240 _0095_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_251_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1248_ net255 _0897_ _0879_ _0896_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1179_ RF.regs\[1\]\[20\] _0862_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ clknet_leaf_24_clk _0194_ _0018_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1038 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2151_ _0005_ net133 _0774_ _0779_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__a31o_1
XFILLER_0_280_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1102_ _0810_ MEM_WB.wb_alu_result\[17\] VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2082_ _0763_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__inv_2
XFILLER_0_233_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1935_ _0746_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1866_ _0620_ _0659_ _0678_ _0679_ _0682_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__a311o_1
XFILLER_0_128_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1797_ _0595_ _0596_ _0610_ _0616_ _0617_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__a311o_1
XFILLER_0_12_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2349_ clknet_leaf_15_clk net344 _0147_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_233_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1720_ _0543_ _0544_ _0545_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__a21oi_4
XFILLER_0_182_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1651_ _0420_ _0454_ _0457_ _0475_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__and4_1
XFILLER_0_184_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold108 ID_EX.ex_rs_data\[6\] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold119 _0237_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1582_ _0331_ _1020_ _1066_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__and3b_1
XFILLER_0_46_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2203_ _0748_ net128 _0773_ _0807_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2134_ _0747_ net104 _0953_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2065_ _0762_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1918_ _0732_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1849_ ID_EX.ex_rt_data\[27\] net123 _0563_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_1211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1703_ _0527_ _0528_ _0529_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1634_ _0390_ _0461_ _0463_ _1042_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1565_ _0395_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__xor2_4
XFILLER_0_26_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1496_ _0321_ _0332_ _0325_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__nor3_1
XFILLER_0_225_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2117_ _0767_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2048_ _0760_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__inv_2
XFILLER_0_230_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1012 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_236_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1350_ _0950_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_263_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1281_ net93 _0913_ net377 VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_274_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_194_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1617_ _0403_ _0429_ _0446_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__a21o_1
XFILLER_0_258_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2597_ net11 VGND VGND VPWR VPWR _2597_/X sky130_fd_sc_hd__buf_2
XFILLER_0_125_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1548_ _0343_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_227_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1479_ _1021_ _0316_ _1034_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_281_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcpu_top_149 VGND VGND VPWR VPWR cpu_top_149/HI dbg_instr[7] sky130_fd_sc_hd__conb_1
XFILLER_0_46_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_249_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2520_ net68 VGND VGND VPWR VPWR _2520_/X sky130_fd_sc_hd__buf_2
XFILLER_0_183_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1402_ net73 VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2382_ clknet_leaf_17_clk net204 _0180_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1333_ net99 _0901_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__or2_1
XFILLER_0_276_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1264_ net375 _0852_ _0002_ _0844_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1195_ net299 _0865_ _0877_ _0868_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_9355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_232_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1951_ _0751_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1882_ _0352_ _0697_ _0698_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2503_ net91 VGND VGND VPWR VPWR _2503_/X sky130_fd_sc_hd__buf_2
XFILLER_0_45_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2365_ clknet_leaf_26_clk net51 _0163_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_224_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_282_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1316_ net76 _0931_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_276_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2296_ clknet_leaf_4_clk net244 _0094_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_263_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1247_ net284 _0897_ _0877_ _0896_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_194_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1178_ net273 _0865_ _0867_ _0868_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_20 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_192_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2150_ net374 _0769_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__and2_1
XFILLER_0_245_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1101_ _0825_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_4
XFILLER_0_89_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2081_ _0763_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__inv_2
XFILLER_0_219_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_232_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1934_ net1 VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1865_ _0670_ _0680_ _0681_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1796_ _0606_ _0615_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2417_ clknet_leaf_18_clk _0314_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2348_ clknet_leaf_15_clk net391 _0146_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2279_ clknet_leaf_10_clk net297 _0077_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_251_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1650_ _0454_ _0457_ _0475_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold109 _0251_ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1581_ _1049_ _1067_ _0331_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__nor3_1
XFILLER_0_61_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_240_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2202_ net363 _0768_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2133_ _0768_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__buf_2
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2064_ _0762_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1917_ _0352_ _0730_ _0731_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__and3_1
XFILLER_0_161_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1848_ _0383_ net60 VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1779_ _0601_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_4
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_264_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1702_ _0497_ _0511_ _0483_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__and3b_1
XFILLER_0_42_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1633_ _0353_ _0462_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1564_ _1011_ _0396_ _0397_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__o21a_2
XFILLER_0_199_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1495_ _1058_ _0319_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_265_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_234_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2116_ _0746_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2047_ _0760_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1020 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_241_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1280_ net389 _0914_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_831 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1616_ _0403_ _0429_ _0446_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__nand3_1
X_2596_ net10 VGND VGND VPWR VPWR _2596_/X sky130_fd_sc_hd__buf_2
XFILLER_0_26_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1547_ net105 ID_EX.ex_rs_data\[10\] _0381_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1478_ _0315_ net70 VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_250_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_245_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1401_ _0994_ _0997_ _0993_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2381_ clknet_leaf_16_clk net214 _0179_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1332_ net100 _0941_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1263_ _0899_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__buf_1
XFILLER_0_120_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1194_ RF.regs\[1\]\[13\] _0875_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__and2_1
XFILLER_0_189_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2579_ net2 VGND VGND VPWR VPWR _2579_/X sky130_fd_sc_hd__buf_2
XFILLER_0_285_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_227_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1950_ _0749_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1881_ _0683_ _0696_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__nand2_2
XFILLER_0_126_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2502_ net90 VGND VGND VPWR VPWR _2502_/X sky130_fd_sc_hd__buf_2
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2364_ clknet_leaf_1_clk net332 _0162_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1315_ net75 _0903_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2295_ clknet_leaf_3_clk net228 _0093_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1246_ net229 _0897_ _0876_ _0896_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1177_ _0844_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_10 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_21 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_284_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_9197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1100_ _0810_ MEM_WB.wb_alu_result\[18\] VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__and2b_1
XFILLER_0_206_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2080_ _0763_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1933_ net97 VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1864_ _0670_ _0680_ _0654_ _0675_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__o211a_1
XFILLER_0_245_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1795_ _0606_ _0615_ _0611_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2416_ clknet_leaf_18_clk _0313_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_274_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2347_ clknet_leaf_18_clk net395 _0145_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2278_ clknet_leaf_10_clk net283 _0076_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1229_ net298 _0890_ _0858_ _0894_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_212_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_270_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_249_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1580_ _0409_ _0412_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_277_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2201_ _0748_ net127 _0773_ _0806_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2132_ _0746_ _0953_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2063_ _0762_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1916_ _0694_ _0698_ _0710_ _0712_ _0728_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__a311o_1
XFILLER_0_127_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1847_ _0621_ _0639_ _0653_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__and3b_2
XFILLER_0_114_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1778_ _0352_ _0599_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_207_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_268_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1701_ _0495_ _0509_ _0510_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__o21a_1
XFILLER_0_121_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1632_ ID_EX.ex_rt_data\[15\] net110 _0373_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_285_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1563_ _1011_ _0391_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1494_ _1064_ _0326_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_254_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2115_ _0766_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__inv_2
XFILLER_0_234_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2046_ _0760_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_256_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1032 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1055 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1615_ _0390_ _0443_ _0445_ _1042_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__a211o_1
XFILLER_0_125_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2595_ net9 VGND VGND VPWR VPWR _2595_/X sky130_fd_sc_hd__buf_2
XFILLER_0_239_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1546_ _1012_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__buf_4
XFILLER_0_238_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1477_ net73 VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_281_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2029_ _0759_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_247_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1400_ _0980_ _0998_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__nor2_4
XFILLER_0_27_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2380_ clknet_leaf_8_clk EX_MEM.rd_in\[1\] _0178_ VGND VGND VPWR VPWR EX_MEM.mem_rd\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_283_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1331_ net99 _0901_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_276_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1262_ ID.CU.ctrl_alusrc _0849_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__and2_1
XFILLER_0_263_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1193_ net261 _0865_ _0876_ _0868_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_203_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_273_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2578_ net128 VGND VGND VPWR VPWR _2578_/X sky130_fd_sc_hd__buf_2
XFILLER_0_168_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1529_ _0362_ _0363_ _0359_ _0360_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_226_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_282_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1880_ _0683_ _0696_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_261_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1097 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2501_ net89 VGND VGND VPWR VPWR _2501_/X sky130_fd_sc_hd__buf_2
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2363_ clknet_leaf_1_clk net392 _0161_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1314_ _0930_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2294_ clknet_leaf_5_clk net264 _0092_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1245_ _0846_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1176_ RF.regs\[1\]\[21\] _0862_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__and2_1
XFILLER_0_189_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_11 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_9110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_266_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1932_ _0744_ _0745_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__nor2_8
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1863_ _0673_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1794_ _0609_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2415_ clknet_leaf_8_clk _0312_ VGND VGND VPWR VPWR RF.regs\[1\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_271_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2346_ clknet_leaf_18_clk net378 _0144_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2277_ clknet_leaf_9_clk _0250_ _0075_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1228_ net235 _0890_ _0857_ _0894_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1159_ net276 _0853_ _0857_ _0855_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__a22o_1
XFILLER_0_181_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_240_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ net338 _0768_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__and2_1
XTAP_7593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_266_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2131_ _0749_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2062_ _0762_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1915_ _0728_ _0729_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__nand2_1
XFILLER_0_267_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_245_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_249_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1846_ _0664_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_115_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1777_ _0596_ _0598_ _0595_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_974 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2329_ clknet_leaf_8_clk net16 _0127_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dfrtp_4
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1056 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_279_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_235_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1066 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_264_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1700_ _0525_ _0526_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1631_ _0343_ net47 VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1562_ net106 ID_EX.ex_rs_data\[11\] _1012_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _0330_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_4
XFILLER_0_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_280_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2114_ _0766_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__inv_2
XFILLER_0_207_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2045_ _0760_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1829_ _0647_ _0648_ _0969_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_257_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1044 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_246_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1067 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1614_ _0353_ _0444_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2594_ net8 VGND VGND VPWR VPWR _2594_/X sky130_fd_sc_hd__buf_2
XFILLER_0_112_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1545_ _0954_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1476_ ID_EX.ex_rt_data\[7\] net133 _1003_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2028_ _0753_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_268_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1330_ _0940_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_258_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1261_ net313 _0852_ _0893_ HAZ.if_id_rt\[0\] VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1192_ RF.regs\[1\]\[14\] _0875_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2577_ net127 VGND VGND VPWR VPWR _2577_/X sky130_fd_sc_hd__buf_2
XFILLER_0_220_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1528_ _0359_ _0360_ _0362_ _0363_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1459_ net73 net69 VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__or2b_1
XFILLER_0_255_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_9347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_268_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1053 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2500_ net88 VGND VGND VPWR VPWR _2500_/X sky130_fd_sc_hd__buf_2
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2362_ clknet_leaf_12_clk net385 _0160_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1313_ _0904_ _0929_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__and2b_1
XFILLER_0_276_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2293_ clknet_leaf_1_clk net274 _0091_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_263_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1244_ net223 _0895_ _0874_ _0896_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__a22o_1
XFILLER_0_223_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1175_ net263 _0865_ _0866_ _0855_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_12 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput130 net130 VGND VGND VPWR VPWR dbg_wb[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_9111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1931_ _0726_ _0731_ _0743_ _0980_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__a31o_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1862_ _0658_ _0660_ _0674_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__and3_1
XFILLER_0_284_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1793_ _0595_ _0597_ _0610_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2414_ clknet_leaf_11_clk _0311_ VGND VGND VPWR VPWR RF.regs\[1\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2345_ clknet_leaf_18_clk net398 _0143_ VGND VGND VPWR VPWR MEM_WB.wb_memtoreg sky130_fd_sc_hd__dfrtp_1
XFILLER_0_271_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2276_ clknet_leaf_15_clk net327 _0074_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_237_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1227_ net330 _0890_ _0856_ _0894_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__a22o_1
XFILLER_0_237_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1158_ RF.regs\[1\]\[29\] _0004_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1089_ _0819_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_4
XFILLER_0_176_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_283_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2130_ _0749_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__inv_2
XFILLER_0_252_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_266_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2061_ _0753_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__buf_4
XFILLER_0_261_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1914_ _0694_ _0698_ _0710_ _0712_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1845_ _0352_ _0662_ _0663_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1776_ _0595_ _0596_ _0598_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__or3_1
XFILLER_0_163_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_256_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_986 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_272_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2328_ clknet_leaf_3_clk net15 _0126_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dfrtp_4
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2259_ clknet_leaf_0_clk net291 _0057_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1068 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_267_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_270_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1630_ _0454_ _0456_ _0458_ _0460_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__o31a_4
XFILLER_0_281_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1561_ _0377_ _0394_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_238_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1492_ _0969_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__and2_1
XFILLER_0_254_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_254_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2113_ _0766_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__inv_2
XFILLER_0_280_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2044_ _0760_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__inv_2
XFILLER_0_234_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1828_ _0620_ _0632_ _0630_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__a21o_1
XFILLER_0_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap140 net14 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__buf_4
X_1759_ _0343_ net55 VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_257_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1613_ ID_EX.ex_rt_data\[14\] net109 _0373_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2593_ net7 VGND VGND VPWR VPWR _2593_/X sky130_fd_sc_hd__buf_2
XFILLER_0_10_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1544_ _0377_ _0378_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__or2_4
XFILLER_0_199_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1475_ _1065_ _1068_ _1069_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__a21oi_2
XFILLER_0_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2027_ _0758_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1260_ ID_EX.ex_rt_data\[1\] _0852_ _0892_ HAZ.if_id_rt\[0\] VGND VGND VPWR VPWR
+ _0214_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1191_ _0849_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__buf_2
XTAP_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2576_ net125 VGND VGND VPWR VPWR _2576_/X sky130_fd_sc_hd__buf_2
XFILLER_0_112_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1527_ _1011_ _0354_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1458_ ID_EX.ex_rt_data\[6\] net132 _1003_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1389_ _0983_ _0985_ _0987_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_241_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2361_ clknet_leaf_27_clk net370 _0159_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1312_ net76 net75 _0903_ net77 VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2292_ clknet_leaf_1_clk net254 _0090_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1243_ net237 _0895_ _0873_ _0896_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a22o_1
XFILLER_0_237_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1174_ RF.regs\[1\]\[22\] _0862_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_13 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput120 net120 VGND VGND VPWR VPWR dbg_wb[24] sky130_fd_sc_hd__clkbuf_4
Xoutput131 net131 VGND VGND VPWR VPWR dbg_wb[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2559_ net107 VGND VGND VPWR VPWR _2559_/X sky130_fd_sc_hd__buf_2
XFILLER_0_80_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_266_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_214_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1930_ _0726_ net180 _0743_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_139_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1861_ _0658_ _0674_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_245_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1792_ net183 _0612_ _0613_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__a21oi_4
XFILLER_0_25_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2413_ clknet_leaf_6_clk _0310_ VGND VGND VPWR VPWR RF.regs\[1\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2344_ clknet_leaf_8_clk _0280_ _0142_ VGND VGND VPWR VPWR FU.id_ex_rs\[0\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2275_ clknet_leaf_16_clk net318 _0073_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_263_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1226_ net294 _0890_ _0854_ _0894_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__a22o_1
XFILLER_0_233_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1157_ net307 _0853_ _0856_ _0855_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1088_ _0810_ MEM_WB.wb_alu_result\[24\] VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1025 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1069 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_266_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2060_ _0761_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__inv_2
XFILLER_0_221_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1913_ _0726_ _0727_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1844_ _0658_ _0661_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1775_ _0561_ _0597_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_269_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_272_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2327_ clknet_leaf_26_clk net14 _0125_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dfrtp_4
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2258_ clknet_leaf_0_clk net260 _0056_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_224_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1209_ net296 _0878_ _0885_ _0881_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__a22o_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2189_ _0748_ net120 _0773_ _0800_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__a31o_1
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_250_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_246_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1560_ _0390_ _0391_ _0393_ _1042_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__a211o_2
XFILLER_0_2_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1491_ _0326_ _0328_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_266_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2112_ _0766_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__inv_2
XFILLER_0_207_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2043_ _0760_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__inv_2
XFILLER_0_221_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1827_ _0645_ _0646_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1758_ _0581_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_4
XFILLER_0_111_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1689_ net113 _0373_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_198_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_898 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_250_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_196_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_246_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1612_ _0343_ net46 VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__nand2_1
XFILLER_0_285_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2592_ net6 VGND VGND VPWR VPWR _2592_/X sky130_fd_sc_hd__buf_2
XFILLER_0_160_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1543_ _0321_ _0358_ _0376_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1474_ _1065_ _1068_ _0969_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_254_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2026_ _0758_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_232_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1190_ net309 _0865_ _0874_ _0868_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__a22o_1
XTAP_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2575_ net124 VGND VGND VPWR VPWR _2575_/X sky130_fd_sc_hd__buf_2
XFILLER_0_239_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1526_ _1011_ _0361_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1457_ _1050_ _1051_ _1052_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__o21a_4
XFILLER_0_215_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1388_ _0964_ _0986_ EX_MEM.ex_memread VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__a21o_1
XFILLER_0_236_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2009_ _0757_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_282_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_230_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_268_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2360_ clknet_leaf_1_clk net393 _0158_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1311_ _0928_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2291_ clknet_leaf_0_clk net246 _0089_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1242_ net241 _0895_ _0872_ _0896_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__a22o_1
XFILLER_0_223_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1173_ _0852_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_256_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_14 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput110 net110 VGND VGND VPWR VPWR dbg_wb[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput121 net121 VGND VGND VPWR VPWR dbg_wb[25] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput132 net132 VGND VGND VPWR VPWR dbg_wb[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2558_ net106 VGND VGND VPWR VPWR _2558_/X sky130_fd_sc_hd__buf_2
XFILLER_0_112_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1509_ _0341_ _0345_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__nor2_1
XFILLER_0_273_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2489_ net77 VGND VGND VPWR VPWR _2489_/X sky130_fd_sc_hd__buf_2
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_266_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1860_ _0674_ _0676_ _0677_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__a21oi_4
XFILLER_0_210_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1791_ _0610_ _0612_ _0969_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2412_ clknet_leaf_7_clk _0309_ VGND VGND VPWR VPWR RF.regs\[1\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2343_ clknet_leaf_9_clk _0279_ _0141_ VGND VGND VPWR VPWR ID.CU.ctrl_alusrc sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2274_ clknet_leaf_16_clk net336 _0072_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1225_ HAZ.if_id_rt\[0\] VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1156_ RF.regs\[1\]\[30\] _0004_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1087_ _0818_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_244_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1989_ _0755_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1912_ _0721_ _0725_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__or2_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1843_ _0658_ _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1774_ _0556_ _0575_ _0576_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_142_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_6_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2326_ clknet_leaf_1_clk net12 _0124_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_209_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2257_ clknet_leaf_0_clk net242 _0055_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_280_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1208_ RF.regs\[1\]\[7\] _0875_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__and2_1
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2188_ net357 _0795_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__and2_1
XFILLER_0_192_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1139_ _0844_ HAZ.if_id_rt\[0\] FU.id_ex_rt\[0\] EX_MEM.ex_memread VGND VGND VPWR
+ VPWR _0845_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _1065_ _1068_ _0327_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__o21a_1
XTAP_8072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2111_ _0766_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2042_ _0760_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1826_ _0640_ _0641_ _0644_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1757_ _0969_ _0580_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__and2_1
XFILLER_0_269_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1688_ ID_EX.ex_rt_data\[18\] net198 VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__nand2_1
XFILLER_0_256_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2309_ clknet_leaf_14_clk net24 _0107_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dfrtp_4
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1611_ _0442_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_4
XFILLER_0_41_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2591_ net141 VGND VGND VPWR VPWR _2591_/X sky130_fd_sc_hd__buf_2
XFILLER_0_23_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1542_ _0321_ _0358_ _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__and3_2
XFILLER_0_23_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1473_ _1020_ _1066_ _1067_ _1049_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_103_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2025_ _0758_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_888 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1809_ _0626_ _0629_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold220 net59 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_271_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_263_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_235_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_250_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_242_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2574_ net123 VGND VGND VPWR VPWR _2574_/X sky130_fd_sc_hd__buf_2
XFILLER_0_125_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1525_ net135 ID_EX.ex_rs_data\[9\] net195 VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1456_ _1050_ _1051_ _0980_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_254_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1387_ net73 net63 VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_207_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2008_ _0757_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_218_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1310_ _0926_ _0927_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__and2_1
XFILLER_0_282_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2290_ clknet_leaf_0_clk net289 _0088_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_236_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1241_ net259 _0895_ _0871_ _0896_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1172_ net227 _0853_ _0864_ _0855_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__a22o_1
XFILLER_0_251_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_15 net142 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput100 net100 VGND VGND VPWR VPWR dbg_pc[6] sky130_fd_sc_hd__clkbuf_4
Xoutput111 net111 VGND VGND VPWR VPWR dbg_wb[16] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_203_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput122 net122 VGND VGND VPWR VPWR dbg_wb[26] sky130_fd_sc_hd__clkbuf_4
Xoutput133 net133 VGND VGND VPWR VPWR dbg_wb[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2557_ net105 VGND VGND VPWR VPWR _2557_/X sky130_fd_sc_hd__buf_2
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1508_ _0954_ _0342_ _0344_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2488_ net76 VGND VGND VPWR VPWR _2488_/X sky130_fd_sc_hd__buf_2
XFILLER_0_255_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_270_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1439_ ID_EX.ex_rt_data\[5\] net196 VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_281_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1790_ _0611_ _0600_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2411_ clknet_leaf_5_clk _0308_ VGND VGND VPWR VPWR RF.regs\[1\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_284_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2342_ clknet_leaf_16_clk _0278_ _0140_ VGND VGND VPWR VPWR HAZ.if_id_rs\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_237_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2273_ clknet_leaf_16_clk net322 _0071_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1224_ net275 _0890_ _0893_ _0844_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1155_ net301 _0853_ _0854_ _0855_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1086_ _0811_ MEM_WB.wb_alu_result\[25\] VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1988_ _0755_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2609_ net25 VGND VGND VPWR VPWR _2609_/X sky130_fd_sc_hd__buf_2
XFILLER_0_140_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_8232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1911_ _0721_ _0725_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__nand2_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1842_ _0620_ _0659_ _0660_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1773_ _0578_ _0575_ _0576_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__o21a_1
XFILLER_0_269_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2325_ clknet_leaf_26_clk net11 _0123_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dfrtp_4
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2256_ clknet_leaf_6_clk net238 _0054_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1207_ net249 _0878_ _0884_ _0881_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__a22o_1
XFILLER_0_224_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2187_ _0788_ net119 _0773_ _0799_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__a31o_1
XFILLER_0_178_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1138_ HAZ.if_id_rs\[0\] VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__buf_2
XFILLER_0_149_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_268_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_672 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_266_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2110_ _0766_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2041_ _0760_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1825_ _0640_ _0641_ _0644_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1756_ _0577_ _0579_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1687_ _0514_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ clknet_leaf_18_clk net13 _0106_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dfrtp_4
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2239_ clknet_leaf_9_clk net174 _0037_ VGND VGND VPWR VPWR ID_EX.ex_aluop\[0\] sky130_fd_sc_hd__dfstp_4
XFILLER_0_280_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1015 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1610_ _0352_ _0440_ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2590_ net4 VGND VGND VPWR VPWR _2590_/X sky130_fd_sc_hd__buf_2
XFILLER_0_23_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1541_ _0983_ _0372_ _0374_ _0375_ _1034_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__a311o_1
XFILLER_0_142_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1472_ _1030_ _1048_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_254_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2024_ _0758_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1808_ _0383_ net57 _0573_ _0628_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold210 net90 VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold221 net52 VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__dlygate4sd3_1
X_1739_ _0373_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_229_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_258_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2573_ net122 VGND VGND VPWR VPWR _2573_/X sky130_fd_sc_hd__buf_2
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1524_ _0321_ _0340_ _0357_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1455_ _1020_ _1032_ _1030_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1386_ _0984_ _0841_ net400 VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2007_ _0757_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_9307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1240_ net290 _0895_ _0870_ _0896_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1171_ RF.regs\[1\]\[23\] _0862_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__and2_1
XFILLER_0_204_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_16 net142 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_261_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput101 net101 VGND VGND VPWR VPWR dbg_pc[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput112 net112 VGND VGND VPWR VPWR dbg_wb[17] sky130_fd_sc_hd__clkbuf_4
Xoutput123 net123 VGND VGND VPWR VPWR dbg_wb[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput134 net134 VGND VGND VPWR VPWR dbg_wb[8] sky130_fd_sc_hd__clkbuf_4
X_2556_ net135 VGND VGND VPWR VPWR _2556_/X sky130_fd_sc_hd__buf_2
XFILLER_0_112_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1507_ _0343_ net71 _0951_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__and3_1
XFILLER_0_255_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2487_ net75 VGND VGND VPWR VPWR _2487_/X sky130_fd_sc_hd__buf_2
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1438_ EX_MEM.ex_memread VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_254_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1369_ _0967_ _0968_ _0969_ VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__o21a_4
XFILLER_0_39_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1020 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_232_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2410_ clknet_leaf_7_clk _0307_ VGND VGND VPWR VPWR RF.regs\[1\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2341_ clknet_leaf_16_clk _0277_ _0139_ VGND VGND VPWR VPWR HAZ.if_id_rt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_283_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2272_ clknet_leaf_17_clk _0245_ _0070_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_236_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1223_ RF.regs\[1\]\[0\] _0849_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__and2_1
XFILLER_0_272_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1154_ _0844_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1085_ _0817_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_220_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1987_ _0755_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_283_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2608_ net23 VGND VGND VPWR VPWR _2608_/X sky130_fd_sc_hd__buf_2
XFILLER_0_140_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2539_ net57 VGND VGND VPWR VPWR _2539_/X sky130_fd_sc_hd__buf_2
XFILLER_0_41_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_254_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_946 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_268_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1910_ _0724_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1841_ _0630_ _0645_ _0646_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_38_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_284_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1772_ _0590_ _0594_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2324_ clknet_leaf_26_clk net10 _0122_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dfrtp_4
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2255_ clknet_leaf_0_clk net224 _0053_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1206_ RF.regs\[1\]\[8\] _0875_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__and2_1
X_2186_ net368 _0795_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1137_ _0843_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_152_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2040_ _0760_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__inv_2
XFILLER_0_221_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1824_ _0573_ _0642_ _0643_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1755_ _0556_ _0561_ _0578_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_41_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1686_ _0352_ _0512_ _0513_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_245_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2307_ clknet_leaf_17_clk net2 _0105_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfrtp_4
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2238_ clknet_leaf_9_clk net376 _0036_ VGND VGND VPWR VPWR ID_EX.ex_imm\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_224_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2169_ net356 _0782_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__and2_1
XFILLER_0_240_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_281_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_868 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1540_ _1000_ net42 _0983_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1471_ _1032_ _1050_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2023_ _0758_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__inv_2
XFILLER_0_261_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1807_ _0380_ _0627_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold200 RF.regs\[1\]\[7\] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold211 net48 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold222 net56 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__dlygate4sd3_1
X_1738_ _0556_ _0561_ _0562_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__a21oi_2
XFILLER_0_142_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1669_ _0483_ _0497_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__xor2_2
XFILLER_0_111_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2572_ net121 VGND VGND VPWR VPWR _2572_/X sky130_fd_sc_hd__buf_2
XFILLER_0_124_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1523_ _0321_ _0358_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1454_ _1048_ _1049_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__nor2_1
XFILLER_0_254_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1385_ ID_EX.ex_rt_data\[2\] VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__inv_2
XFILLER_0_207_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_253_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2006_ _0753_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__buf_4
XFILLER_0_171_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2239__174 VGND VGND VPWR VPWR net174 _2239__174/LO sky130_fd_sc_hd__conb_1
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ net243 _0853_ _0863_ _0855_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_218_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_254_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_17 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput102 net102 VGND VGND VPWR VPWR dbg_pc[8] sky130_fd_sc_hd__clkbuf_4
Xoutput113 net113 VGND VGND VPWR VPWR dbg_wb[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput124 net124 VGND VGND VPWR VPWR dbg_wb[28] sky130_fd_sc_hd__buf_2
XFILLER_0_203_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput135 net135 VGND VGND VPWR VPWR dbg_wb[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2555_ net134 VGND VGND VPWR VPWR _2555_/X sky130_fd_sc_hd__buf_2
XFILLER_0_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_259_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1506_ _1000_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2486_ net74 VGND VGND VPWR VPWR _2486_/X sky130_fd_sc_hd__buf_2
XFILLER_0_254_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1437_ net192 _1032_ _1033_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__o21a_4
XFILLER_0_255_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_270_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1368_ ID_EX.ex_aluop\[0\] VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_173_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1299_ net83 _0906_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__nor2_1
XFILLER_0_214_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_271_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_204_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2340_ clknet_leaf_8_clk net203 _0138_ VGND VGND VPWR VPWR EX_MEM.mem_regwrite sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2271_ clknet_leaf_9_clk net295 _0069_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_229_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1222_ net321 _0890_ _0892_ _0844_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_252_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1153_ RF.regs\[1\]\[31\] _0004_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__and2_1
XFILLER_0_220_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1084_ _0811_ MEM_WB.wb_alu_result\[26\] VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1986_ _0755_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_9_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2607_ net22 VGND VGND VPWR VPWR _2607_/X sky130_fd_sc_hd__buf_2
XFILLER_0_247_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2538_ net56 VGND VGND VPWR VPWR _2538_/X sky130_fd_sc_hd__buf_2
XFILLER_0_122_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_254_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_249_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1080 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_266_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_273_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_260_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1840_ _0632_ _0647_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1771_ _0491_ _0592_ _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_108_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2323_ clknet_leaf_25_clk net9 _0121_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dfrtp_4
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2254_ clknet_leaf_6_clk net230 _0052_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1205_ net319 _0878_ _0883_ _0881_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2185_ _0788_ net118 _0786_ _0798_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1136_ MEM_WB.wb_memtoreg MEM_WB.wb_alu_result\[0\] VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1969_ _0752_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_233_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_268_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_279_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1823_ _0573_ _0635_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1754_ _0551_ _0555_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1685_ _0495_ _0499_ _0511_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ clknet_leaf_8_clk _0004_ _0104_ VGND VGND VPWR VPWR EX_MEM.ex_regwrite sky130_fd_sc_hd__dfrtp_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2237_ clknet_leaf_23_clk _0211_ _0035_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_252_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2168_ _0788_ net109 _0786_ _0789_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__a31o_1
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1119_ _0834_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_4
XFILLER_0_36_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2099_ _0765_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__inv_2
XFILLER_0_230_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_247_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1470_ _1064_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__inv_2
XFILLER_0_266_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2022_ _0758_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__inv_2
XFILLER_0_221_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1050 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_253_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1806_ net120 ID_EX.ex_rs_data\[24\] _0591_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold201 ID_EX.ex_imm\[12\] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold212 net57 VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__dlygate4sd3_1
X_1737_ _0556_ _0561_ _0969_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__o21ai_1
Xhold223 net65 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1668_ _0495_ _0496_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__or2_2
XFILLER_0_121_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1599_ _0403_ _0408_ _0428_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__a21o_1
XFILLER_0_238_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2571_ net120 VGND VGND VPWR VPWR _2571_/X sky130_fd_sc_hd__buf_2
XFILLER_0_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1522_ _0340_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1453_ _1046_ _1047_ _1041_ _1044_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_284_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1384_ _0982_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__buf_4
XFILLER_0_222_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2005_ _0756_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_872 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_254_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_18 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_248_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput103 net103 VGND VGND VPWR VPWR dbg_pc[9] sky130_fd_sc_hd__buf_2
XFILLER_0_101_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput114 net114 VGND VGND VPWR VPWR dbg_wb[19] sky130_fd_sc_hd__clkbuf_4
X_2554_ net133 VGND VGND VPWR VPWR _2554_/X sky130_fd_sc_hd__buf_2
Xoutput125 net125 VGND VGND VPWR VPWR dbg_wb[29] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput136 net179 VGND VGND VPWR VPWR dbg_wb_rd[0] sky130_fd_sc_hd__buf_2
XFILLER_0_140_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1505_ net134 ID_EX.ex_rs_data\[8\] _1012_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_267_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2485_ net103 VGND VGND VPWR VPWR _2485_/X sky130_fd_sc_hd__buf_2
XFILLER_0_103_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1436_ _1020_ _1032_ _0980_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_254_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_270_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1367_ _0966_ _0957_ _0959_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__and3_1
XFILLER_0_270_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1298_ net84 _0907_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__xor2_1
XFILLER_0_222_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2270_ clknet_leaf_9_clk net331 _0068_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_256_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1221_ RF.regs\[1\]\[1\] _0849_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__and2_1
XFILLER_0_236_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1152_ _0852_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1083_ _0816_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1985_ _0755_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2606_ net21 VGND VGND VPWR VPWR _2606_/X sky130_fd_sc_hd__buf_2
XFILLER_0_28_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2537_ net55 VGND VGND VPWR VPWR _2537_/X sky130_fd_sc_hd__buf_2
XFILLER_0_268_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1419_ _1014_ _1015_ _1010_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__a21o_1
XFILLER_0_215_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2399_ clknet_leaf_0_clk _0296_ VGND VGND VPWR VPWR RF.regs\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1770_ _0491_ _0582_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2322_ clknet_leaf_26_clk net8 _0120_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dfrtp_4
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2253_ clknet_leaf_6_clk net285 _0051_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1204_ RF.regs\[1\]\[9\] _0875_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2184_ net360 _0795_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__and2_1
XFILLER_0_251_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1135_ _0842_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_6
XFILLER_0_178_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1968_ _0752_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1899_ _0352_ _0713_ _0714_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1822_ net121 ID_EX.ex_rs_data\[25\] _0591_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1753_ _0575_ _0576_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__and2b_1
XFILLER_0_53_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1684_ _0495_ _0499_ _0511_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ clknet_leaf_9_clk _0002_ _0103_ VGND VGND VPWR VPWR EX_MEM.ex_memread sky130_fd_sc_hd__dfrtp_4
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2236_ clknet_leaf_23_clk _0210_ _0034_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_212_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_234_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2167_ net359 _0782_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__and2_1
XFILLER_0_221_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1118_ _0809_ MEM_WB.wb_alu_result\[9\] VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__and2b_1
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2098_ _0765_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_241_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_250_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2021_ _0758_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__inv_2
XFILLER_0_206_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1062 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_253_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1805_ _0621_ _0625_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1736_ _0483_ _0557_ _0559_ _0560_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__a211oi_2
Xhold202 _0212_ VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold213 net45 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold224 net73 VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_269_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1667_ _0490_ _0494_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__and2_1
XFILLER_0_284_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1598_ _0403_ _0429_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2219_ clknet_leaf_21_clk _0193_ _0017_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_197_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2570_ net119 VGND VGND VPWR VPWR _2570_/X sky130_fd_sc_hd__buf_2
XFILLER_0_129_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1521_ _0353_ _0354_ _0356_ _1034_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__a211o_1
XFILLER_0_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1452_ _1041_ _1044_ _1046_ _1047_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__o211a_1
XFILLER_0_266_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1383_ FU.id_ex_rt\[0\] _0949_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__nand2_1
XFILLER_0_282_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_222_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2004_ _0756_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__inv_2
XFILLER_0_270_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1719_ _0543_ _0544_ _0969_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_269_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_245_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_19 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput104 net104 VGND VGND VPWR VPWR dbg_wb[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_242_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput115 net115 VGND VGND VPWR VPWR dbg_wb[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2553_ net132 VGND VGND VPWR VPWR _2553_/X sky130_fd_sc_hd__buf_2
Xoutput126 net126 VGND VGND VPWR VPWR dbg_wb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_100_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput137 net175 VGND VGND VPWR VPWR dbg_wb_rd[1] sky130_fd_sc_hd__buf_2
XFILLER_0_267_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1504_ net191 _0340_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2484_ net102 VGND VGND VPWR VPWR _2484_/X sky130_fd_sc_hd__buf_2
XFILLER_0_107_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1435_ _1030_ _1031_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1366_ _0957_ _0959_ _0966_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_282_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1297_ _0908_ _0921_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_246_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_220_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_248_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1220_ net335 _0890_ _0891_ _0881_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1151_ _0846_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_251_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1082_ _0811_ MEM_WB.wb_alu_result\[27\] VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__and2b_1
XFILLER_0_220_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1984_ _0753_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__buf_4
XFILLER_0_51_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2605_ net20 VGND VGND VPWR VPWR _2605_/X sky130_fd_sc_hd__buf_2
XFILLER_0_261_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2536_ net54 VGND VGND VPWR VPWR _2536_/X sky130_fd_sc_hd__buf_2
XFILLER_0_228_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1418_ _1010_ _1014_ _1015_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__and3_1
XFILLER_0_254_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2398_ clknet_leaf_5_clk _0295_ VGND VGND VPWR VPWR RF.regs\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_270_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1349_ FU.id_ex_rs\[0\] _0949_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_233_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_240_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1042 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_283_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2321_ clknet_leaf_1_clk net7 _0119_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_283_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2252_ clknet_leaf_11_clk net256 _0050_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_280_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1203_ net315 _0878_ _0882_ _0881_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2183_ _0788_ net117 _0786_ _0797_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__a31o_1
XFILLER_0_252_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1134_ MEM_WB.wb_memtoreg MEM_WB.wb_alu_result\[1\] VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__or2_1
XFILLER_0_215_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1967_ _0752_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1898_ _0711_ _0712_ _0694_ _0698_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_47_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2519_ net67 VGND VGND VPWR VPWR _2519_/X sky130_fd_sc_hd__buf_2
XFILLER_0_41_1036 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_268_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_285_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1821_ _0621_ _0625_ _0638_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_38_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1752_ _0572_ _0574_ _0569_ _0570_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__a211o_1
XFILLER_0_147_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1683_ _0509_ _0510_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_267_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2304_ clknet_leaf_8_clk _0003_ _0102_ VGND VGND VPWR VPWR ID_EX.ex_regdst sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ clknet_leaf_23_clk _0209_ _0033_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_213_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2166_ _0748_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1117_ _0833_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2097_ _0765_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__inv_2
XFILLER_0_234_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_278_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2020_ _0758_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__inv_2
XFILLER_0_250_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1074 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1804_ _0585_ _0624_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__and2b_1
XFILLER_0_182_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1735_ _0495_ _0509_ _0510_ _0527_ _0543_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold203 net95 VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold214 net42 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_257_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold225 net53 VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1666_ _0490_ _0494_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1597_ _0408_ _0428_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__and2_4
XFILLER_0_102_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_237_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2218_ clknet_leaf_14_clk _0192_ _0016_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_252_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2149_ _0005_ net132 _0774_ _0778_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1520_ _1021_ _0355_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1451_ _1011_ _1037_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_267_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1382_ _0966_ _0973_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__nand2_1
XFILLER_0_248_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_250_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2003_ _0756_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_231_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_277_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1718_ _0525_ _0531_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__nand2_2
XFILLER_0_203_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1649_ _0478_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_0_284_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_260_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_269_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_248_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1022 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_259_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput105 net105 VGND VGND VPWR VPWR dbg_wb[10] sky130_fd_sc_hd__clkbuf_4
X_2552_ net131 VGND VGND VPWR VPWR _2552_/X sky130_fd_sc_hd__buf_2
XFILLER_0_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput116 net116 VGND VGND VPWR VPWR dbg_wb[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput127 net127 VGND VGND VPWR VPWR dbg_wb[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput138 net178 VGND VGND VPWR VPWR dbg_wb_we sky130_fd_sc_hd__clkbuf_4
X_1503_ _0338_ _0339_ _1034_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__a21o_1
XFILLER_0_267_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2483_ net101 VGND VGND VPWR VPWR _2483_/X sky130_fd_sc_hd__buf_2
XFILLER_0_282_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1434_ _1026_ _1029_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_281_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1365_ _0961_ _0965_ _0958_ _0964_ EX_MEM.ex_memread VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__a221o_2
XFILLER_0_128_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_235_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1296_ net84 _0907_ net85 VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_250_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_277_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_248_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1150_ _0851_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_232_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1081_ _0815_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1983_ _0754_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2604_ net19 VGND VGND VPWR VPWR _2604_/X sky130_fd_sc_hd__buf_2
XFILLER_0_140_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2535_ net53 VGND VGND VPWR VPWR _2535_/X sky130_fd_sc_hd__buf_2
XFILLER_0_109_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1417_ _1011_ _1001_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2397_ clknet_leaf_6_clk _0294_ VGND VGND VPWR VPWR RF.regs\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_254_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1348_ EX_MEM.mem_rd\[1\] EX_MEM.mem_regwrite EX_MEM.mem_rd\[0\] VGND VGND VPWR VPWR
+ _0949_ sky130_fd_sc_hd__and3b_1
XFILLER_0_93_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1279_ net95 net93 _0913_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2320_ clknet_leaf_25_clk net6 _0118_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dfrtp_4
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2251_ clknet_leaf_11_clk net222 _0049_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1202_ RF.regs\[1\]\[10\] _0875_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2182_ net365 _0795_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__and2_1
XFILLER_0_217_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1133_ _0841_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__inv_4
XFILLER_0_251_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1966_ _0752_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__inv_2
XFILLER_0_267_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1897_ _0694_ _0698_ _0711_ _0712_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__a211o_1
XFILLER_0_70_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2518_ net66 VGND VGND VPWR VPWR _2518_/X sky130_fd_sc_hd__buf_2
XFILLER_0_59_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1820_ _0621_ _0639_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_167_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1751_ _0569_ _0570_ _0572_ _0574_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1682_ _0505_ _0508_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__or2_4
XFILLER_0_123_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ clknet_leaf_8_clk net302 _0101_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_267_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2234_ clknet_leaf_23_clk _0208_ _0032_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dfrtp_4
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2165_ _0005_ net108 _0786_ _0787_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1116_ _0810_ MEM_WB.wb_alu_result\[10\] VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2096_ _0765_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__inv_2
XFILLER_0_230_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1949_ _0750_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_280_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_250_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_250_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_203_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1803_ _0383_ net57 _0546_ _0623_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1734_ _0539_ _0542_ _0558_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold204 net41 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 net96 VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1665_ _0491_ _0492_ _0493_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_284_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1596_ _0353_ _0425_ _0427_ _1034_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__a211o_1
XFILLER_0_258_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2217_ clknet_leaf_14_clk _0191_ _0015_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2148_ net364 _0769_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2079_ _0763_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__inv_2
XFILLER_0_269_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1450_ ID_EX.ex_rs_data\[5\] _1012_ _1045_ _0951_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__a211o_1
XFILLER_0_266_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1381_ ID_EX.ex_aluop\[0\] VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__inv_6
XFILLER_0_282_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2002_ _0756_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1717_ _0539_ _0542_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__xor2_4
XFILLER_0_44_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1648_ _0352_ _0476_ _0477_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1579_ _0315_ _0406_ _0380_ _0411_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__o31a_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer30 _0960_ VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_269_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1034 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2551_ net130 VGND VGND VPWR VPWR _2551_/X sky130_fd_sc_hd__buf_2
XFILLER_0_281_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput106 net106 VGND VGND VPWR VPWR dbg_wb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_224_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput117 net117 VGND VGND VPWR VPWR dbg_wb[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput128 net128 VGND VGND VPWR VPWR dbg_wb[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1502_ _0983_ _0315_ net71 VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__or3b_1
XFILLER_0_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2482_ net100 VGND VGND VPWR VPWR _2482_/X sky130_fd_sc_hd__buf_2
XFILLER_0_267_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1433_ _1026_ _1029_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__and2_1
XFILLER_0_227_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1364_ ID_EX.ex_rt_data\[0\] _0962_ _0964_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_281_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1295_ _0909_ _0920_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_235_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_270_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_246_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_272_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_248_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1080_ _0811_ MEM_WB.wb_alu_result\[28\] VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__and2b_1
XFILLER_0_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1982_ _0754_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2603_ net18 VGND VGND VPWR VPWR _2603_/X sky130_fd_sc_hd__buf_2
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2534_ net51 VGND VGND VPWR VPWR _2534_/X sky130_fd_sc_hd__buf_2
XFILLER_0_140_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1416_ _1011_ _1013_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__or2_1
XFILLER_0_283_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2396_ clknet_leaf_11_clk _0293_ VGND VGND VPWR VPWR RF.regs\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_242_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1347_ _0948_ VGND VGND VPWR VPWR EX_MEM.rd_in\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_251_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1278_ net92 _0912_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_266_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_271_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ clknet_leaf_10_clk net312 _0048_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1201_ net265 _0878_ _0880_ _0881_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_236_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2181_ _0788_ net116 _0786_ _0796_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1132_ _0809_ MEM_WB.wb_alu_result\[2\] VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__nor2_2
XFILLER_0_75_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_267_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1965_ _0752_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1896_ _0708_ _0709_ _0706_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2517_ net63 VGND VGND VPWR VPWR _2517_/X sky130_fd_sc_hd__buf_2
XFILLER_0_267_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2379_ clknet_leaf_16_clk EX_MEM.rd_in\[0\] _0177_ VGND VGND VPWR VPWR EX_MEM.mem_rd\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_242_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1750_ _0573_ _0565_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_249_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1681_ _0505_ _0508_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2302_ clknet_leaf_9_clk net308 _0100_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2233_ clknet_leaf_23_clk _0207_ _0031_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dfrtp_4
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2164_ net342 _0782_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_273_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1115_ _0832_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_4
XFILLER_0_221_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2095_ _0765_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1948_ _0750_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1879_ _0694_ _0695_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__and2_1
XFILLER_0_241_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1802_ ID_EX.ex_rt_data\[24\] _0563_ _0622_ _0983_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1733_ _0539_ _0542_ _0525_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold205 EX_MEM.ex_memread VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold216 ID_EX.ex_regdst VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1664_ _0491_ _0484_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1595_ _0353_ _0426_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2216_ clknet_leaf_21_clk _0190_ _0014_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_252_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_234_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2147_ net210 _0769_ _0777_ _0774_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2078_ _0763_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1380_ net187 net190 _0979_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__a21boi_4
XFILLER_0_281_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2001_ _0756_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_270_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_203_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1716_ _0491_ _0540_ _0541_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_124_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_258_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1647_ _0452_ _0459_ _0475_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__or3_1
XFILLER_0_258_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1578_ _0380_ _0410_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_258_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer20 net193 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__buf_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer31 _0402_ VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_269_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_206_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_263_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1046 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2550_ net129 VGND VGND VPWR VPWR _2550_/X sky130_fd_sc_hd__buf_2
XFILLER_0_106_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput107 net107 VGND VGND VPWR VPWR dbg_wb[12] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_259_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput118 net118 VGND VGND VPWR VPWR dbg_wb[22] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput129 net129 VGND VGND VPWR VPWR dbg_wb[3] sky130_fd_sc_hd__buf_2
X_1501_ _0983_ _0337_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2481_ net99 VGND VGND VPWR VPWR _2481_/X sky130_fd_sc_hd__buf_2
XFILLER_0_220_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_259_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1432_ _0951_ _1023_ _1028_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_266_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1363_ _0963_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__buf_2
XFILLER_0_282_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1294_ net86 _0908_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__nor2_1
XFILLER_0_235_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1029 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_268_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_248_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_219_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1981_ _0754_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__inv_2
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2602_ net17 VGND VGND VPWR VPWR _2602_/X sky130_fd_sc_hd__buf_2
XFILLER_0_148_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2533_ net50 VGND VGND VPWR VPWR _2533_/X sky130_fd_sc_hd__buf_2
XFILLER_0_267_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1415_ net129 ID_EX.ex_rs_data\[3\] _1012_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_243_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2395_ clknet_leaf_11_clk _0292_ VGND VGND VPWR VPWR RF.regs\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1346_ FU.id_ex_rs\[0\] net390 VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1277_ net91 net90 _0911_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_285_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1200_ _0844_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_280_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2180_ net351 _0795_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1131_ _0840_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__buf_4
XFILLER_0_233_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1964_ _0752_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_808 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1895_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_259_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_243_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2516_ net52 VGND VGND VPWR VPWR _2516_/X sky130_fd_sc_hd__buf_2
XFILLER_0_45_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_227_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_243_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2378_ clknet_leaf_8_clk net212 _0176_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1329_ _0902_ _0939_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__and2b_1
XFILLER_0_270_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1018 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1680_ _0491_ _0506_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__o21a_1
XFILLER_0_52_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_8581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_267_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_249_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2301_ clknet_leaf_7_clk net277 _0099_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2232_ clknet_leaf_23_clk _0206_ _0030_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dfrtp_4
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2163_ _0953_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1114_ _0810_ MEM_WB.wb_alu_result\[11\] VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__and2b_1
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2094_ _0746_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_178_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1947_ _0750_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1878_ _0690_ _0693_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_257_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1801_ net120 net199 VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1732_ _0497_ _0511_ _0527_ _0543_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__and4b_1
XFILLER_0_170_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold206 net81 VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__dlygate4sd3_1
X_1663_ net111 ID_EX.ex_rs_data\[16\] _0381_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__mux2_1
Xhold217 net63 VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_262_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_9090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_285_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_278_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1594_ ID_EX.ex_rt_data\[13\] net108 net182 VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_240_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2215_ clknet_leaf_21_clk _0189_ _0013_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dfrtp_4
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2146_ _0749_ _0838_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_178_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2077_ _0763_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2000_ _0756_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_690 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1715_ _0491_ _0533_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_258_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1646_ _0452_ _0459_ _0475_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1577_ net107 ID_EX.ex_rs_data\[12\] _0381_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer10 _0402_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__buf_6
XFILLER_0_69_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer21 _0955_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2129_ _0749_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_269_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1500_ ID_EX.ex_rt_data\[8\] net134 _1003_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput108 net108 VGND VGND VPWR VPWR dbg_wb[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput119 net119 VGND VGND VPWR VPWR dbg_wb[23] sky130_fd_sc_hd__buf_2
XFILLER_0_51_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2480_ net98 VGND VGND VPWR VPWR _2480_/X sky130_fd_sc_hd__buf_2
XFILLER_0_224_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1431_ _0839_ net194 _1027_ _0954_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1362_ EX_MEM.mem_rd\[1\] EX_MEM.mem_regwrite FU.id_ex_rt\[0\] EX_MEM.mem_rd\[0\]
+ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__and4b_1
XFILLER_0_120_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput90 net90 VGND VGND VPWR VPWR dbg_pc[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_247_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_235_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1293_ net87 _0909_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__xor2_1
XFILLER_0_250_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1629_ _0980_ _0459_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_285_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_260_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_248_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1980_ _0754_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2601_ net16 VGND VGND VPWR VPWR _2601_/X sky130_fd_sc_hd__buf_2
Xrebuffer1 net137 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2532_ net49 VGND VGND VPWR VPWR _2532_/X sky130_fd_sc_hd__buf_2
XFILLER_0_12_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1414_ _0955_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2394_ clknet_leaf_6_clk _0291_ VGND VGND VPWR VPWR RF.regs\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_259_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1345_ _0947_ VGND VGND VPWR VPWR EX_MEM.rd_in\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_282_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1276_ net89 _0910_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1130_ MEM_WB.wb_memtoreg MEM_WB.wb_alu_result\[3\] VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__and2b_1
XFILLER_0_256_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_267_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1963_ _0752_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__inv_2
XFILLER_0_267_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1894_ _0706_ _0708_ _0709_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__or3_4
XFILLER_0_128_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2515_ net41 VGND VGND VPWR VPWR _2515_/X sky130_fd_sc_hd__buf_2
XFILLER_0_278_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2377_ clknet_leaf_3_clk net397 _0175_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_236_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1328_ net100 net99 _0901_ net101 VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__a31o_1
XFILLER_0_169_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1259_ net339 _0852_ _0891_ _0898_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_231_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_242_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_9261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_8571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2300_ clknet_leaf_8_clk net287 _0098_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ clknet_leaf_23_clk _0205_ _0029_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dfrtp_4
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2162_ _0005_ net107 _0774_ _0785_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__a31o_1
XFILLER_0_178_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1113_ _0831_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_4
XFILLER_0_24_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2093_ _0764_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_267_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1946_ _0750_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1877_ _0690_ _0693_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1800_ _0538_ _0568_ _0587_ _0605_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__or4b_4
XFILLER_0_143_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1731_ _0551_ _0555_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_198_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1662_ _0432_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__buf_4
XFILLER_0_83_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold207 net69 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold218 net49 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1593_ _1000_ net45 VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ clknet_leaf_14_clk _0188_ _0012_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dfrtp_4
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2145_ net209 _0769_ _0776_ _0774_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__a22o_1
XFILLER_0_252_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2076_ _0763_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1929_ _0739_ _0742_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_280_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold90 _0267_ VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_264_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1714_ net114 ID_EX.ex_rs_data\[19\] _0381_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_258_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1645_ _0472_ _0474_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1576_ _0403_ _0408_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__xor2_1
XFILLER_0_272_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_226_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer11 net401 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer22 _0962_ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2128_ _0749_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__inv_2
XFILLER_0_174_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1040 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2059_ _0761_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__inv_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_241_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_276_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_250_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput109 net109 VGND VGND VPWR VPWR dbg_wb[14] sky130_fd_sc_hd__buf_2
XFILLER_0_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1430_ ID_EX.ex_rs_data\[4\] net194 VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1361_ net137 net176 FU.id_ex_rt\[0\] net136 VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_248_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput80 net80 VGND VGND VPWR VPWR dbg_pc[16] sky130_fd_sc_hd__buf_2
Xoutput91 net91 VGND VGND VPWR VPWR dbg_pc[27] sky130_fd_sc_hd__buf_2
XFILLER_0_281_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1292_ _0910_ _0919_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__nor2_1
XFILLER_0_272_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1628_ _0456_ _0458_ _0454_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1559_ _0353_ _0392_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_202_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2600_ net15 VGND VGND VPWR VPWR _2600_/X sky130_fd_sc_hd__buf_2
XFILLER_0_148_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer2 net138 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__buf_1
XFILLER_0_10_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2531_ net48 VGND VGND VPWR VPWR _2531_/X sky130_fd_sc_hd__buf_2
XFILLER_0_45_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1413_ _0951_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_259_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2393_ clknet_leaf_9_clk _0290_ VGND VGND VPWR VPWR RF.regs\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1344_ ID_EX.ex_regdst FU.id_ex_rt\[0\] VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__and2b_1
XFILLER_0_276_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1275_ net88 net87 _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__and3_2
XFILLER_0_250_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_233_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_267_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_248_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1962_ _0752_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1893_ FU.id_ex_rs\[0\] _0949_ _0700_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2514_ net39 VGND VGND VPWR VPWR _2514_/X sky130_fd_sc_hd__buf_2
XFILLER_0_60_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2376_ clknet_leaf_12_clk net64 _0174_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_255_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1327_ _0938_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1258_ net303 _0852_ _0889_ _0898_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1189_ RF.regs\[1\]\[15\] _0862_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ clknet_leaf_19_clk _0204_ _0028_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_264_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2161_ net341 _0782_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1112_ _0809_ MEM_WB.wb_alu_result\[12\] VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2092_ _0764_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__inv_2
XFILLER_0_191_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1945_ _0750_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__inv_2
XFILLER_0_267_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1876_ _0315_ _0687_ _0380_ _0692_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__o31a_1
XFILLER_0_128_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2359_ clknet_leaf_25_clk net387 _0157_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_249_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1730_ _0554_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1661_ _0488_ _0489_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__nor2_1
Xhold208 net62 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 net46 VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1592_ _0409_ _0412_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2213_ clknet_leaf_14_clk _0187_ _0011_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dfrtp_4
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2144_ _0749_ _0839_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2075_ _0763_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1928_ _0573_ _0740_ _0741_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1036 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1859_ _0674_ _0676_ _0969_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_285_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 _0265_ VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_264_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold91 ID_EX.ex_rs_data\[11\] VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_251_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1713_ _0520_ _0536_ _0538_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__o21a_2
XFILLER_0_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1644_ _0473_ _0471_ _0468_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__or3b_4
XFILLER_0_83_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1575_ _1034_ _0405_ _0407_ _1039_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__o31a_1
XFILLER_0_26_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer12 _1025_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer23 net196 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__buf_1
XFILLER_0_94_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2127_ _0749_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__inv_2
XFILLER_0_221_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2058_ _0761_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__inv_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_280_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_249_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput2 net2 VGND VGND VPWR VPWR dbg_alu[0] sky130_fd_sc_hd__buf_2
XFILLER_0_220_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1360_ net104 _0960_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__nand2_1
Xoutput70 net70 VGND VGND VPWR VPWR dbg_mem_addr[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput81 net81 VGND VGND VPWR VPWR dbg_pc[17] sky130_fd_sc_hd__clkbuf_4
Xoutput92 net92 VGND VGND VPWR VPWR dbg_pc[28] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_247_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1291_ net87 _0909_ net88 VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_194_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_203_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1627_ _0417_ _0420_ _0457_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__o21a_1
XFILLER_0_258_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1558_ ID_EX.ex_rt_data\[11\] net106 _0373_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_258_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_226_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1489_ _1058_ _1059_ _1063_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_241_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_245_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer3 net176 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__buf_1
XFILLER_0_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2530_ net47 VGND VGND VPWR VPWR _2530_/X sky130_fd_sc_hd__buf_2
XFILLER_0_122_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1412_ _1006_ net201 VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2392_ clknet_leaf_10_clk _0289_ VGND VGND VPWR VPWR RF.regs\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1343_ net208 _0853_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_237_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1274_ net86 _0908_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__and2_1
XFILLER_0_235_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1043 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_215_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_262_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_205_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1961_ _0749_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__buf_6
XFILLER_0_16_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_248_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1892_ _0573_ _0707_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2513_ net39 VGND VGND VPWR VPWR _2513_/X sky130_fd_sc_hd__buf_2
XFILLER_0_243_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_5_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_259_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2375_ clknet_leaf_25_clk net382 _0173_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1326_ _0936_ _0937_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_235_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1257_ net328 _0852_ _0888_ _0898_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__a22o_1
XFILLER_0_250_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1188_ net280 _0865_ _0873_ _0868_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_231_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_248_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_8573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_221_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2160_ _0005_ net106 _0774_ _0784_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__a31o_1
XFILLER_0_261_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1111_ _0830_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_4
XFILLER_0_233_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2091_ _0764_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_232_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_267_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1944_ _0750_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1875_ _0380_ _0691_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2358_ clknet_leaf_12_clk net366 _0156_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1309_ net78 _0904_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__or2_1
XTAP_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2289_ clknet_leaf_0_clk net248 _0087_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_251_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_947 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_249_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1660_ _0403_ _0466_ _0487_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold209 net67 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_9071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1591_ _0413_ _0421_ _0423_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_260_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2212_ clknet_leaf_13_clk _0186_ _0010_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_265_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2143_ _0005_ net129 _0774_ _0775_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__a31o_1
XFILLER_0_234_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2074_ _0763_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1927_ _0573_ _0733_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1858_ _0654_ _0675_ _0663_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_142_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1789_ _0588_ _0589_ _0594_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_275_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold70 _0269_ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold81 ID_EX.ex_rt_data\[12\] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold92 _0256_ VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1712_ net184 _0466_ _0537_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__nand3_4
XFILLER_0_26_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 _0810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1643_ net185 _0466_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1574_ _0315_ _0406_ _1021_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__o21a_1
XFILLER_0_238_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2126_ _0767_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__inv_2
Xrebuffer13 _0967_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_1
XFILLER_0_136_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer24 net197 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_1
XFILLER_0_156_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2057_ _0761_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__inv_2
XFILLER_0_178_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1041 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_275_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_223_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_265_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_239_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput3 net3 VGND VGND VPWR VPWR dbg_alu[10] sky130_fd_sc_hd__buf_2
XFILLER_0_122_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_254_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput60 net60 VGND VGND VPWR VPWR dbg_mem_addr[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_247_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput71 net71 VGND VGND VPWR VPWR dbg_mem_addr[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_263_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput82 net82 VGND VGND VPWR VPWR dbg_pc[18] sky130_fd_sc_hd__buf_2
XFILLER_0_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput93 net93 VGND VGND VPWR VPWR dbg_pc[29] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_207_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1290_ _0911_ _0918_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_216_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1626_ _0438_ _0413_ _0436_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_83_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_285_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1557_ _0343_ net43 VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_273_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_266_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1488_ _0322_ _0325_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2109_ _0766_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_241_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_241_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer4 net177 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__buf_4
XFILLER_0_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1411_ _1008_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__buf_6
XFILLER_0_121_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2391_ clknet_leaf_10_clk _0288_ VGND VGND VPWR VPWR RF.regs\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1342_ _0946_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1273_ net85 net84 _0907_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__and3_1
XFILLER_0_257_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_250_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1055 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1609_ _0424_ _0422_ _0439_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_258_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2589_ net3 VGND VGND VPWR VPWR _2589_/X sky130_fd_sc_hd__buf_2
XFILLER_0_274_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_247_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1960_ _0751_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__inv_2
XFILLER_0_189_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_248_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1891_ net125 ID_EX.ex_rs_data\[29\] _0591_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2512_ net39 VGND VGND VPWR VPWR _2512_/X sky130_fd_sc_hd__buf_2
XFILLER_0_122_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2374_ clknet_leaf_7_clk net61 _0172_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_242_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1325_ net102 _0902_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_282_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1256_ net323 _0897_ _0887_ _0898_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1187_ RF.regs\[1\]\[16\] _0862_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_226_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_9297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_224_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_217_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1110_ _0809_ MEM_WB.wb_alu_result\[13\] VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__and2b_1
XFILLER_0_156_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2090_ _0764_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__inv_2
XFILLER_0_233_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_956 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1943_ _0750_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1874_ net124 ID_EX.ex_rs_data\[28\] _0591_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_243_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2357_ clknet_leaf_12_clk net369 _0155_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1308_ net79 _0926_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2288_ clknet_leaf_0_clk net281 _0086_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_212_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1239_ net217 _0895_ _0869_ _0896_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__a22o_1
XFILLER_0_212_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_222_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_959 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire141 net5 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__buf_4
XFILLER_0_80_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ _0980_ _0422_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2211_ clknet_leaf_13_clk _0185_ _0009_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_256_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_280_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2142_ net367 _0769_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__and2_1
XFILLER_0_179_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2073_ _0763_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1926_ net128 ID_EX.ex_rs_data\[31\] _0591_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1857_ _0657_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1788_ _0606_ _0609_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_204_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2409_ clknet_leaf_5_clk _0306_ VGND VGND VPWR VPWR RF.regs\[1\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_274_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold60 _0235_ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold71 ID_EX.ex_rs_data\[19\] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold82 _0225_ VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold93 ID_EX.ex_rs_data\[12\] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_268_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_213_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1711_ _0504_ _0519_ _0536_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_2 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1642_ _0467_ _0468_ _0471_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_112_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1573_ net44 VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer14 _0731_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
X_2125_ _0767_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__inv_2
XFILLER_0_234_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer25 net197 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_179_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2056_ _0761_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_251_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_838 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_228_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1909_ _0315_ _0718_ _0380_ _0723_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__o31a_1
XFILLER_0_60_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_283_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput4 net4 VGND VGND VPWR VPWR dbg_alu[11] sky130_fd_sc_hd__buf_2
XFILLER_0_202_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput50 net50 VGND VGND VPWR VPWR dbg_mem_addr[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput61 net61 VGND VGND VPWR VPWR dbg_mem_addr[28] sky130_fd_sc_hd__clkbuf_4
Xoutput72 net72 VGND VGND VPWR VPWR dbg_mem_addr[9] sky130_fd_sc_hd__buf_2
XFILLER_0_275_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput83 net83 VGND VGND VPWR VPWR dbg_pc[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput94 net94 VGND VGND VPWR VPWR dbg_pc[2] sky130_fd_sc_hd__buf_2
XFILLER_0_208_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_262_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1025 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_186_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_207_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1625_ _0455_ _0436_ _0438_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_78_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1556_ _0353_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1487_ _0323_ _0324_ _0954_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_281_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2108_ _0766_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2039_ _0753_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_254_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_252_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer5 net136 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_210_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1410_ _0966_ _0973_ _1007_ _1005_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__and4_1
XFILLER_0_62_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2390_ clknet_leaf_9_clk _0287_ VGND VGND VPWR VPWR RF.regs\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_236_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1341_ HAZ.if_id_rt\[0\] _0852_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__or2_1
XFILLER_0_247_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_237_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1272_ net83 _0906_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__and2_1
XFILLER_0_263_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_270_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1040 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_270_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1068 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_248_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1067 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_190_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1608_ _0424_ _0422_ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_273_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2588_ net33 VGND VGND VPWR VPWR _2588_/X sky130_fd_sc_hd__buf_2
XFILLER_0_239_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_220_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1539_ net105 _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_226_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_282_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_227_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_199_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_231_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_208_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold190 RF.regs\[1\]\[6\] VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_232_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1890_ _0704_ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2511_ net36 VGND VGND VPWR VPWR _2511_/X sky130_fd_sc_hd__buf_2
XFILLER_0_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2373_ clknet_leaf_27_clk net60 _0171_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1324_ net103 _0936_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_270_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_208_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_223_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1255_ net251 _0897_ _0886_ _0898_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_250_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1186_ net247 _0865_ _0872_ _0868_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__a22o_1
XFILLER_0_231_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_270_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_231_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_231_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_214_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_252_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_206_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1942_ _0750_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__inv_2
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1873_ _0684_ _0689_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__xor2_1
XFILLER_0_160_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_226_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2356_ clknet_leaf_6_clk net388 _0154_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1307_ net78 _0904_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2287_ clknet_leaf_6_clk net310 _0085_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_251_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1238_ net225 _0895_ _0867_ _0896_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_237_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1169_ RF.regs\[1\]\[24\] _0862_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_285_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_261_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_274_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_255_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_203_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_284_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1060 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire142 net30 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__buf_4
XFILLER_0_81_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_269_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2210_ clknet_leaf_14_clk _0184_ _0008_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dfrtp_4
XTAP_7693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2141_ _0773_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_280_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2072_ _0753_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_233_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1925_ _0737_ _0738_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__nor2_1
XFILLER_0_267_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_695 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1856_ _0670_ _0673_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_167_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1787_ _0491_ _0607_ _0608_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_278_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2408_ clknet_leaf_5_clk _0305_ VGND VGND VPWR VPWR RF.regs\[1\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_243_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_283_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2339_ clknet_leaf_17_clk net379 _0137_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dfrtp_4
XTAP_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_246_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold50 _0228_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold61 ID_EX.ex_rt_data\[29\] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold72 _0264_ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold83 ID_EX.ex_rs_data\[27\] VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_243_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold94 _0257_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_264_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1710_ _0390_ _0533_ _0535_ _1042_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1641_ _0432_ _0469_ _0470_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__o21a_1
XANTENNA_3 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1572_ _0353_ _0404_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2124_ _0767_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__inv_2
XFILLER_0_238_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_222_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer15 _0978_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_1
Xrebuffer26 _0999_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_171_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_233_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2055_ _0761_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_212_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_282_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1908_ _0380_ _0722_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1839_ _0654_ _0657_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_274_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_246_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput5 net141 VGND VGND VPWR VPWR dbg_alu[12] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput40 net40 VGND VGND VPWR VPWR dbg_instr[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_222_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput51 net51 VGND VGND VPWR VPWR dbg_mem_addr[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput62 net62 VGND VGND VPWR VPWR dbg_mem_addr[29] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput73 net73 VGND VGND VPWR VPWR dbg_memread sky130_fd_sc_hd__clkbuf_4
Xoutput84 net84 VGND VGND VPWR VPWR dbg_pc[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_207_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput95 net95 VGND VGND VPWR VPWR dbg_pc[30] sky130_fd_sc_hd__clkbuf_4
XTAP_6063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_262_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1624_ _0409_ _0412_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__or2_1
XFILLER_0_257_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1555_ _0389_ VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_4
XFILLER_0_26_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1486_ net133 ID_EX.ex_rs_data\[7\] _1012_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2107_ _0766_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_19_clk clknet_1_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2038_ _0759_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_276_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_244_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer6 net188 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_63_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_239_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_241_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1340_ net94 _0852_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_208_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_263_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1271_ net82 net81 _0905_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__and3_1
XFILLER_0_262_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1052 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1079 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_clk clknet_1_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_125_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1607_ _0437_ _0438_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2587_ net32 VGND VGND VPWR VPWR _2587_/X sky130_fd_sc_hd__buf_2
XFILLER_0_41_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_273_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1538_ net181 VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__buf_6
XFILLER_0_61_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_220_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1469_ _1060_ _1063_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_227_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_236_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_236_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_175_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_282_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_247_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_8768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold180 RF.regs\[1\]\[27\] VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold191 RF.regs\[1\]\[21\] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_218_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_244_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_260_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_269_1481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_1329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2510_ net35 VGND VGND VPWR VPWR _2510_/X sky130_fd_sc_hd__buf_2
XFILLER_0_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_183_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2372_ clknet_leaf_7_clk net394 _0170_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1323_ net102 _0902_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_264_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_263_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_271_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_276_1485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1254_ net271 _0897_ _0885_ _0898_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1185_ RF.regs\[1\]\[17\] _0862_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_270_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_231_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_231_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_273_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_1661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_226_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_282_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_241_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_1509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_255_1569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_210_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_194_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_266_1621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_1605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_1665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_1649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_9255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_8576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_245_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_273_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_261_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_1609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_219_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_216_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_213_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1941_ _0750_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_210_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_189_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1872_ _0983_ _0685_ _0686_ _0688_ _0585_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__a311o_1
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_245_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_265_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_209_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2355_ clknet_leaf_15_clk net372 _0153_ VGND VGND VPWR VPWR MEM_WB.wb_alu_result\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_271_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_208_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_264_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1306_ _0925_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_223_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2286_ clknet_leaf_6_clk net262 _0084_ VGND VGND VPWR VPWR ID_EX.ex_rs_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_224_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_252_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1237_ HAZ.if_id_rt\[0\] VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_233_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1168_ _0849_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__buf_2
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_250_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1099_ _0824_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__buf_4
XFILLER_0_177_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_176_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_1024 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_244_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_228_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_227_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_216_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_242_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_255_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_214_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_214_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_284_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1072 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_262_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_227_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_184_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_9063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_9096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _0953_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__clkbuf_4
XTAP_6993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_238_1553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2071_ _0762_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__inv_2
XFILLER_0_227_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_1597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_233_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_191_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_232_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_234_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1924_ _0704_ _0720_ _0736_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249_1693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1855_ _0573_ _0671_ _0672_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1786_ _0491_ _0602_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_256_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_269_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_198_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_256_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_200_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2407_ clknet_leaf_5_clk _0304_ VGND VGND VPWR VPWR RF.regs\[1\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_243_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2338_ clknet_leaf_8_clk net26 _0136_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_271_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_1653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_225_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2269_ clknet_leaf_7_clk net236 _0067_ VGND VGND VPWR VPWR ID_EX.ex_rt_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_251_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_224_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217_1637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_252_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_212_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_177_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_285_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_279_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_263_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_275_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_261_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_248_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_219_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_194_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold40 EX_MEM.mem_rd\[0\] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold51 ID_EX.ex_rt_data\[21\] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold62 _0242_ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold73 ID_EX.ex_rs_data\[17\] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold84 _0272_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold95 ID_EX.ex_rt_data\[8\] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_270_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_215_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_1497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_196_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1640_ _1011_ _0461_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_4 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_227_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_269_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1571_ ID_EX.ex_rt_data\[12\] net107 net181 VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_285_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_240_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_284_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_8170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_1465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_238_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_8192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_238_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_7480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_280_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_207_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2123_ _0767_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__inv_2
XFILLER_0_240_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_280_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_233_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_206_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer16 _0978_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__buf_1
XFILLER_0_179_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1061 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer27 _1009_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_1
X_2054_ _0761_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_202_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_267_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_228_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1907_ net127 ID_EX.ex_rs_data\[30\] _0591_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_267_1089 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_245_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_1633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1838_ _0380_ _0655_ _0656_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_128_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182_1677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_248_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1016 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1769_ net118 ID_EX.ex_rs_data\[22\] _0591_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_257_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_204_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_272_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_283_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_218_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_274_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278_1185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_1049 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_217_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_256_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_1101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_252_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_212_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_178_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_211_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_250_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230_1689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_211_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_192_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228_1541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_180_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_267_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_259_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput6 net6 VGND VGND VPWR VPWR dbg_alu[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_266_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput30 net142 VGND VGND VPWR VPWR dbg_alu[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput41 net41 VGND VGND VPWR VPWR dbg_mem_addr[0] sky130_fd_sc_hd__clkbuf_4
Xoutput52 net52 VGND VGND VPWR VPWR dbg_mem_addr[1] sky130_fd_sc_hd__buf_2
XFILLER_0_43_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_222_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_6020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput63 net63 VGND VGND VPWR VPWR dbg_mem_addr[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_275_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_198_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput74 net74 VGND VGND VPWR VPWR dbg_pc[10] sky130_fd_sc_hd__buf_2
XFILLER_0_262_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput85 net85 VGND VGND VPWR VPWR dbg_pc[21] sky130_fd_sc_hd__buf_2
XFILLER_0_207_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput96 net96 VGND VGND VPWR VPWR dbg_pc[31] sky130_fd_sc_hd__buf_2
XFILLER_0_78_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_257_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_235_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257_1269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_1681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_187_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_204_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_230_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_224_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_1397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_268_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_264_1229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_207_1625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1623_ _0452_ _0453_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_239_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_199_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1554_ _0387_ ID_EX.ex_aluop\[0\] _0388_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__and3b_1
XFILLER_0_239_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_201_1213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_240_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_205_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_254_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1485_ _0316_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__inv_2
XFILLER_0_265_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_1257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_275_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_185_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
.ends

